//`timescale 1ns / 1ps
module bitmap_rom_ddct (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire pixel
);

  reg [7:0] mem[2047:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'hc0;
    mem[116] = 8'h1f;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'hfc;
    mem[132] = 8'hff;
    mem[133] = 8'h03;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'hff;
    mem[140] = 8'h1f;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h80;
    mem[147] = 8'hff;
    mem[148] = 8'hff;
    mem[149] = 8'h1f;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h80;
    mem[155] = 8'hff;
    mem[156] = 8'h3f;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'he0;
    mem[163] = 8'hff;
    mem[164] = 8'hff;
    mem[165] = 8'h7f;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'h80;
    mem[171] = 8'hff;
    mem[172] = 8'h3f;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'hf0;
    mem[179] = 8'hff;
    mem[180] = 8'hff;
    mem[181] = 8'hff;
    mem[182] = 8'h01;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'h80;
    mem[187] = 8'hff;
    mem[188] = 8'h3f;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'hfc;
    mem[195] = 8'hff;
    mem[196] = 8'hff;
    mem[197] = 8'hff;
    mem[198] = 8'h03;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'h00;
    mem[202] = 8'h80;
    mem[203] = 8'hff;
    mem[204] = 8'h3f;
    mem[205] = 8'h00;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'hfe;
    mem[211] = 8'hff;
    mem[212] = 8'hff;
    mem[213] = 8'hff;
    mem[214] = 8'h0f;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'h80;
    mem[219] = 8'hff;
    mem[220] = 8'h3f;
    mem[221] = 8'h00;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'hff;
    mem[227] = 8'hff;
    mem[228] = 8'hff;
    mem[229] = 8'hff;
    mem[230] = 8'h1f;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h80;
    mem[235] = 8'hff;
    mem[236] = 8'h3f;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h80;
    mem[242] = 8'hff;
    mem[243] = 8'hff;
    mem[244] = 8'hff;
    mem[245] = 8'hff;
    mem[246] = 8'h3f;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'h80;
    mem[251] = 8'hff;
    mem[252] = 8'h3f;
    mem[253] = 8'h00;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'hc0;
    mem[258] = 8'hff;
    mem[259] = 8'hff;
    mem[260] = 8'hff;
    mem[261] = 8'hff;
    mem[262] = 8'h7f;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'h80;
    mem[267] = 8'hff;
    mem[268] = 8'h3f;
    mem[269] = 8'h00;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'he0;
    mem[274] = 8'hff;
    mem[275] = 8'hff;
    mem[276] = 8'hff;
    mem[277] = 8'hff;
    mem[278] = 8'h7f;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h80;
    mem[283] = 8'hff;
    mem[284] = 8'h3f;
    mem[285] = 8'h00;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'he0;
    mem[290] = 8'hff;
    mem[291] = 8'hff;
    mem[292] = 8'hff;
    mem[293] = 8'hff;
    mem[294] = 8'hff;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h80;
    mem[299] = 8'hff;
    mem[300] = 8'h3f;
    mem[301] = 8'h00;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'hf0;
    mem[306] = 8'hff;
    mem[307] = 8'hff;
    mem[308] = 8'hff;
    mem[309] = 8'hff;
    mem[310] = 8'hff;
    mem[311] = 8'h01;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h80;
    mem[315] = 8'hff;
    mem[316] = 8'h3f;
    mem[317] = 8'h00;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'hf8;
    mem[322] = 8'hff;
    mem[323] = 8'hff;
    mem[324] = 8'hff;
    mem[325] = 8'hff;
    mem[326] = 8'hff;
    mem[327] = 8'h01;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'h80;
    mem[331] = 8'hff;
    mem[332] = 8'h3f;
    mem[333] = 8'h00;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'hf8;
    mem[338] = 8'hff;
    mem[339] = 8'hff;
    mem[340] = 8'hff;
    mem[341] = 8'hff;
    mem[342] = 8'hff;
    mem[343] = 8'h03;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h80;
    mem[347] = 8'hff;
    mem[348] = 8'h3f;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'hfc;
    mem[354] = 8'hff;
    mem[355] = 8'hff;
    mem[356] = 8'hff;
    mem[357] = 8'hff;
    mem[358] = 8'hff;
    mem[359] = 8'h03;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h80;
    mem[363] = 8'hff;
    mem[364] = 8'h3f;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'hfc;
    mem[370] = 8'hff;
    mem[371] = 8'hff;
    mem[372] = 8'hff;
    mem[373] = 8'hff;
    mem[374] = 8'hff;
    mem[375] = 8'h07;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h80;
    mem[379] = 8'hff;
    mem[380] = 8'h3f;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'hfc;
    mem[386] = 8'hff;
    mem[387] = 8'hff;
    mem[388] = 8'hff;
    mem[389] = 8'hff;
    mem[390] = 8'hff;
    mem[391] = 8'h07;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h80;
    mem[395] = 8'hff;
    mem[396] = 8'h3f;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'hfe;
    mem[402] = 8'hff;
    mem[403] = 8'hff;
    mem[404] = 8'hff;
    mem[405] = 8'hff;
    mem[406] = 8'hff;
    mem[407] = 8'h0f;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h80;
    mem[411] = 8'hff;
    mem[412] = 8'h3f;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'hfe;
    mem[418] = 8'hff;
    mem[419] = 8'hff;
    mem[420] = 8'hff;
    mem[421] = 8'hff;
    mem[422] = 8'hff;
    mem[423] = 8'h0f;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h80;
    mem[427] = 8'hff;
    mem[428] = 8'h7f;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'hfe;
    mem[434] = 8'hff;
    mem[435] = 8'hff;
    mem[436] = 8'hff;
    mem[437] = 8'hff;
    mem[438] = 8'hff;
    mem[439] = 8'h0f;
    mem[440] = 8'hc0;
    mem[441] = 8'hff;
    mem[442] = 8'hff;
    mem[443] = 8'hff;
    mem[444] = 8'hff;
    mem[445] = 8'hff;
    mem[446] = 8'hff;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'hff;
    mem[450] = 8'hff;
    mem[451] = 8'hff;
    mem[452] = 8'hff;
    mem[453] = 8'hff;
    mem[454] = 8'hff;
    mem[455] = 8'h0f;
    mem[456] = 8'he0;
    mem[457] = 8'hff;
    mem[458] = 8'hff;
    mem[459] = 8'hff;
    mem[460] = 8'hff;
    mem[461] = 8'hff;
    mem[462] = 8'hff;
    mem[463] = 8'h01;
    mem[464] = 8'h00;
    mem[465] = 8'hff;
    mem[466] = 8'hff;
    mem[467] = 8'hff;
    mem[468] = 8'hff;
    mem[469] = 8'hff;
    mem[470] = 8'hff;
    mem[471] = 8'h1f;
    mem[472] = 8'he0;
    mem[473] = 8'hff;
    mem[474] = 8'hff;
    mem[475] = 8'hff;
    mem[476] = 8'hff;
    mem[477] = 8'hff;
    mem[478] = 8'hff;
    mem[479] = 8'h01;
    mem[480] = 8'h00;
    mem[481] = 8'hff;
    mem[482] = 8'hff;
    mem[483] = 8'hff;
    mem[484] = 8'hff;
    mem[485] = 8'hff;
    mem[486] = 8'hff;
    mem[487] = 8'h1f;
    mem[488] = 8'he0;
    mem[489] = 8'hff;
    mem[490] = 8'hff;
    mem[491] = 8'hff;
    mem[492] = 8'hff;
    mem[493] = 8'hff;
    mem[494] = 8'hff;
    mem[495] = 8'h01;
    mem[496] = 8'h00;
    mem[497] = 8'hff;
    mem[498] = 8'hff;
    mem[499] = 8'hff;
    mem[500] = 8'hff;
    mem[501] = 8'hff;
    mem[502] = 8'hff;
    mem[503] = 8'h1f;
    mem[504] = 8'he0;
    mem[505] = 8'hff;
    mem[506] = 8'hff;
    mem[507] = 8'hff;
    mem[508] = 8'hff;
    mem[509] = 8'hff;
    mem[510] = 8'hff;
    mem[511] = 8'h01;
    mem[512] = 8'h00;
    mem[513] = 8'hff;
    mem[514] = 8'hff;
    mem[515] = 8'hff;
    mem[516] = 8'hff;
    mem[517] = 8'hff;
    mem[518] = 8'hff;
    mem[519] = 8'h0f;
    mem[520] = 8'he0;
    mem[521] = 8'hff;
    mem[522] = 8'hff;
    mem[523] = 8'hff;
    mem[524] = 8'hff;
    mem[525] = 8'hff;
    mem[526] = 8'hff;
    mem[527] = 8'h01;
    mem[528] = 8'h00;
    mem[529] = 8'hff;
    mem[530] = 8'hff;
    mem[531] = 8'hff;
    mem[532] = 8'hff;
    mem[533] = 8'hff;
    mem[534] = 8'hff;
    mem[535] = 8'h00;
    mem[536] = 8'he0;
    mem[537] = 8'hff;
    mem[538] = 8'hff;
    mem[539] = 8'hff;
    mem[540] = 8'hff;
    mem[541] = 8'hff;
    mem[542] = 8'hff;
    mem[543] = 8'h01;
    mem[544] = 8'h00;
    mem[545] = 8'hff;
    mem[546] = 8'hff;
    mem[547] = 8'hff;
    mem[548] = 8'hff;
    mem[549] = 8'hff;
    mem[550] = 8'h1f;
    mem[551] = 8'h00;
    mem[552] = 8'he0;
    mem[553] = 8'hff;
    mem[554] = 8'hff;
    mem[555] = 8'hff;
    mem[556] = 8'hff;
    mem[557] = 8'hff;
    mem[558] = 8'hff;
    mem[559] = 8'h01;
    mem[560] = 8'h00;
    mem[561] = 8'hff;
    mem[562] = 8'hff;
    mem[563] = 8'hff;
    mem[564] = 8'hff;
    mem[565] = 8'hff;
    mem[566] = 8'h03;
    mem[567] = 8'h00;
    mem[568] = 8'he0;
    mem[569] = 8'hff;
    mem[570] = 8'hff;
    mem[571] = 8'hff;
    mem[572] = 8'hff;
    mem[573] = 8'hff;
    mem[574] = 8'hff;
    mem[575] = 8'h01;
    mem[576] = 8'h00;
    mem[577] = 8'hff;
    mem[578] = 8'hff;
    mem[579] = 8'hff;
    mem[580] = 8'hff;
    mem[581] = 8'hff;
    mem[582] = 8'h01;
    mem[583] = 8'h00;
    mem[584] = 8'he0;
    mem[585] = 8'hff;
    mem[586] = 8'hff;
    mem[587] = 8'hff;
    mem[588] = 8'hff;
    mem[589] = 8'hff;
    mem[590] = 8'hff;
    mem[591] = 8'h01;
    mem[592] = 8'h00;
    mem[593] = 8'hff;
    mem[594] = 8'hff;
    mem[595] = 8'hff;
    mem[596] = 8'hff;
    mem[597] = 8'hff;
    mem[598] = 8'h03;
    mem[599] = 8'h00;
    mem[600] = 8'he0;
    mem[601] = 8'hff;
    mem[602] = 8'hff;
    mem[603] = 8'hff;
    mem[604] = 8'hff;
    mem[605] = 8'hff;
    mem[606] = 8'hff;
    mem[607] = 8'h01;
    mem[608] = 8'h00;
    mem[609] = 8'hfe;
    mem[610] = 8'hff;
    mem[611] = 8'hff;
    mem[612] = 8'hff;
    mem[613] = 8'hff;
    mem[614] = 8'h07;
    mem[615] = 8'h00;
    mem[616] = 8'he0;
    mem[617] = 8'hff;
    mem[618] = 8'hff;
    mem[619] = 8'hff;
    mem[620] = 8'hff;
    mem[621] = 8'hff;
    mem[622] = 8'hff;
    mem[623] = 8'h01;
    mem[624] = 8'h00;
    mem[625] = 8'hfe;
    mem[626] = 8'hff;
    mem[627] = 8'hff;
    mem[628] = 8'hff;
    mem[629] = 8'hff;
    mem[630] = 8'h0f;
    mem[631] = 8'h00;
    mem[632] = 8'he0;
    mem[633] = 8'hff;
    mem[634] = 8'hff;
    mem[635] = 8'hff;
    mem[636] = 8'hff;
    mem[637] = 8'hff;
    mem[638] = 8'hff;
    mem[639] = 8'h01;
    mem[640] = 8'h00;
    mem[641] = 8'hfe;
    mem[642] = 8'hff;
    mem[643] = 8'hff;
    mem[644] = 8'hff;
    mem[645] = 8'hff;
    mem[646] = 8'h3f;
    mem[647] = 8'h00;
    mem[648] = 8'hc0;
    mem[649] = 8'hff;
    mem[650] = 8'hff;
    mem[651] = 8'hff;
    mem[652] = 8'hff;
    mem[653] = 8'hff;
    mem[654] = 8'hff;
    mem[655] = 8'h00;
    mem[656] = 8'h00;
    mem[657] = 8'hfe;
    mem[658] = 8'hff;
    mem[659] = 8'hff;
    mem[660] = 8'hff;
    mem[661] = 8'hff;
    mem[662] = 8'h7f;
    mem[663] = 8'h00;
    mem[664] = 8'h00;
    mem[665] = 8'h00;
    mem[666] = 8'h80;
    mem[667] = 8'hff;
    mem[668] = 8'h7f;
    mem[669] = 8'h00;
    mem[670] = 8'h00;
    mem[671] = 8'h00;
    mem[672] = 8'h00;
    mem[673] = 8'hfc;
    mem[674] = 8'hff;
    mem[675] = 8'hff;
    mem[676] = 8'hff;
    mem[677] = 8'hff;
    mem[678] = 8'hff;
    mem[679] = 8'h00;
    mem[680] = 8'h00;
    mem[681] = 8'h00;
    mem[682] = 8'h80;
    mem[683] = 8'hff;
    mem[684] = 8'h3f;
    mem[685] = 8'h00;
    mem[686] = 8'h00;
    mem[687] = 8'h00;
    mem[688] = 8'h00;
    mem[689] = 8'hfc;
    mem[690] = 8'hff;
    mem[691] = 8'hff;
    mem[692] = 8'hff;
    mem[693] = 8'hff;
    mem[694] = 8'hff;
    mem[695] = 8'h01;
    mem[696] = 8'h00;
    mem[697] = 8'h00;
    mem[698] = 8'h80;
    mem[699] = 8'hff;
    mem[700] = 8'h3f;
    mem[701] = 8'h00;
    mem[702] = 8'h00;
    mem[703] = 8'h00;
    mem[704] = 8'h00;
    mem[705] = 8'hfc;
    mem[706] = 8'hff;
    mem[707] = 8'hff;
    mem[708] = 8'hff;
    mem[709] = 8'hff;
    mem[710] = 8'hff;
    mem[711] = 8'h03;
    mem[712] = 8'h00;
    mem[713] = 8'h00;
    mem[714] = 8'h80;
    mem[715] = 8'hff;
    mem[716] = 8'h3f;
    mem[717] = 8'h00;
    mem[718] = 8'h00;
    mem[719] = 8'h00;
    mem[720] = 8'h00;
    mem[721] = 8'hf8;
    mem[722] = 8'hff;
    mem[723] = 8'hff;
    mem[724] = 8'hff;
    mem[725] = 8'hff;
    mem[726] = 8'hff;
    mem[727] = 8'h03;
    mem[728] = 8'h00;
    mem[729] = 8'h00;
    mem[730] = 8'h80;
    mem[731] = 8'hff;
    mem[732] = 8'h3f;
    mem[733] = 8'h00;
    mem[734] = 8'h00;
    mem[735] = 8'h00;
    mem[736] = 8'h00;
    mem[737] = 8'hf8;
    mem[738] = 8'hff;
    mem[739] = 8'hff;
    mem[740] = 8'hff;
    mem[741] = 8'hff;
    mem[742] = 8'hff;
    mem[743] = 8'h01;
    mem[744] = 8'h00;
    mem[745] = 8'h00;
    mem[746] = 8'h80;
    mem[747] = 8'hff;
    mem[748] = 8'h3f;
    mem[749] = 8'h00;
    mem[750] = 8'h00;
    mem[751] = 8'h00;
    mem[752] = 8'h00;
    mem[753] = 8'hf0;
    mem[754] = 8'hff;
    mem[755] = 8'hff;
    mem[756] = 8'hff;
    mem[757] = 8'hff;
    mem[758] = 8'hff;
    mem[759] = 8'h01;
    mem[760] = 8'h00;
    mem[761] = 8'h00;
    mem[762] = 8'h80;
    mem[763] = 8'hff;
    mem[764] = 8'h3f;
    mem[765] = 8'h00;
    mem[766] = 8'h00;
    mem[767] = 8'h00;
    mem[768] = 8'h00;
    mem[769] = 8'he0;
    mem[770] = 8'hff;
    mem[771] = 8'hff;
    mem[772] = 8'hff;
    mem[773] = 8'hff;
    mem[774] = 8'hff;
    mem[775] = 8'h00;
    mem[776] = 8'h00;
    mem[777] = 8'h00;
    mem[778] = 8'h80;
    mem[779] = 8'hff;
    mem[780] = 8'h3f;
    mem[781] = 8'h00;
    mem[782] = 8'h00;
    mem[783] = 8'h00;
    mem[784] = 8'h00;
    mem[785] = 8'he0;
    mem[786] = 8'hff;
    mem[787] = 8'hff;
    mem[788] = 8'hff;
    mem[789] = 8'hff;
    mem[790] = 8'h7f;
    mem[791] = 8'h00;
    mem[792] = 8'h00;
    mem[793] = 8'h00;
    mem[794] = 8'h80;
    mem[795] = 8'hff;
    mem[796] = 8'h3f;
    mem[797] = 8'h00;
    mem[798] = 8'h00;
    mem[799] = 8'h00;
    mem[800] = 8'h00;
    mem[801] = 8'hc0;
    mem[802] = 8'hff;
    mem[803] = 8'hff;
    mem[804] = 8'hff;
    mem[805] = 8'hff;
    mem[806] = 8'h3f;
    mem[807] = 8'h00;
    mem[808] = 8'h00;
    mem[809] = 8'h00;
    mem[810] = 8'h80;
    mem[811] = 8'hff;
    mem[812] = 8'h3f;
    mem[813] = 8'h00;
    mem[814] = 8'h00;
    mem[815] = 8'h00;
    mem[816] = 8'h00;
    mem[817] = 8'h80;
    mem[818] = 8'hff;
    mem[819] = 8'hff;
    mem[820] = 8'hff;
    mem[821] = 8'hff;
    mem[822] = 8'h1f;
    mem[823] = 8'h00;
    mem[824] = 8'h00;
    mem[825] = 8'h00;
    mem[826] = 8'h80;
    mem[827] = 8'hff;
    mem[828] = 8'h3f;
    mem[829] = 8'h00;
    mem[830] = 8'h00;
    mem[831] = 8'h00;
    mem[832] = 8'h00;
    mem[833] = 8'h00;
    mem[834] = 8'hff;
    mem[835] = 8'hff;
    mem[836] = 8'hff;
    mem[837] = 8'hff;
    mem[838] = 8'h0f;
    mem[839] = 8'h00;
    mem[840] = 8'h00;
    mem[841] = 8'h00;
    mem[842] = 8'h80;
    mem[843] = 8'hff;
    mem[844] = 8'h3f;
    mem[845] = 8'h00;
    mem[846] = 8'h00;
    mem[847] = 8'h00;
    mem[848] = 8'h00;
    mem[849] = 8'h00;
    mem[850] = 8'hfe;
    mem[851] = 8'hff;
    mem[852] = 8'hff;
    mem[853] = 8'hff;
    mem[854] = 8'h07;
    mem[855] = 8'h00;
    mem[856] = 8'h00;
    mem[857] = 8'h00;
    mem[858] = 8'h80;
    mem[859] = 8'hff;
    mem[860] = 8'h3f;
    mem[861] = 8'h00;
    mem[862] = 8'h00;
    mem[863] = 8'h00;
    mem[864] = 8'h00;
    mem[865] = 8'h00;
    mem[866] = 8'hf8;
    mem[867] = 8'hff;
    mem[868] = 8'hff;
    mem[869] = 8'hff;
    mem[870] = 8'h03;
    mem[871] = 8'h00;
    mem[872] = 8'h00;
    mem[873] = 8'h00;
    mem[874] = 8'h80;
    mem[875] = 8'hff;
    mem[876] = 8'h3f;
    mem[877] = 8'h00;
    mem[878] = 8'h00;
    mem[879] = 8'h00;
    mem[880] = 8'h00;
    mem[881] = 8'h00;
    mem[882] = 8'hf0;
    mem[883] = 8'hff;
    mem[884] = 8'hff;
    mem[885] = 8'hff;
    mem[886] = 8'h00;
    mem[887] = 8'h00;
    mem[888] = 8'h00;
    mem[889] = 8'h00;
    mem[890] = 8'h80;
    mem[891] = 8'hff;
    mem[892] = 8'h3f;
    mem[893] = 8'h00;
    mem[894] = 8'h00;
    mem[895] = 8'h00;
    mem[896] = 8'h00;
    mem[897] = 8'h00;
    mem[898] = 8'hc0;
    mem[899] = 8'hff;
    mem[900] = 8'hff;
    mem[901] = 8'h3f;
    mem[902] = 8'h00;
    mem[903] = 8'h00;
    mem[904] = 8'h00;
    mem[905] = 8'h00;
    mem[906] = 8'h80;
    mem[907] = 8'hff;
    mem[908] = 8'h3f;
    mem[909] = 8'h00;
    mem[910] = 8'h00;
    mem[911] = 8'h00;
    mem[912] = 8'h00;
    mem[913] = 8'h00;
    mem[914] = 8'h00;
    mem[915] = 8'hff;
    mem[916] = 8'hff;
    mem[917] = 8'h0f;
    mem[918] = 8'h00;
    mem[919] = 8'h00;
    mem[920] = 8'h00;
    mem[921] = 8'h00;
    mem[922] = 8'h80;
    mem[923] = 8'hff;
    mem[924] = 8'h3f;
    mem[925] = 8'h00;
    mem[926] = 8'h00;
    mem[927] = 8'h00;
    mem[928] = 8'h00;
    mem[929] = 8'h00;
    mem[930] = 8'h00;
    mem[931] = 8'hf8;
    mem[932] = 8'hff;
    mem[933] = 8'h03;
    mem[934] = 8'h00;
    mem[935] = 8'h00;
    mem[936] = 8'h00;
    mem[937] = 8'h00;
    mem[938] = 8'h00;
    mem[939] = 8'hff;
    mem[940] = 8'h1f;
    mem[941] = 8'h00;
    mem[942] = 8'h00;
    mem[943] = 8'h00;
    mem[944] = 8'h00;
    mem[945] = 8'h00;
    mem[946] = 8'h00;
    mem[947] = 8'h00;
    mem[948] = 8'h1f;
    mem[949] = 8'h00;
    mem[950] = 8'h00;
    mem[951] = 8'h00;
    mem[952] = 8'h00;
    mem[953] = 8'h00;
    mem[954] = 8'h00;
    mem[955] = 8'h00;
    mem[956] = 8'h00;
    mem[957] = 8'h00;
    mem[958] = 8'h00;
    mem[959] = 8'h00;
    mem[960] = 8'h00;
    mem[961] = 8'h00;
    mem[962] = 8'h00;
    mem[963] = 8'h00;
    mem[964] = 8'h00;
    mem[965] = 8'h00;
    mem[966] = 8'h00;
    mem[967] = 8'h00;
    mem[968] = 8'h00;
    mem[969] = 8'h00;
    mem[970] = 8'h00;
    mem[971] = 8'h00;
    mem[972] = 8'h00;
    mem[973] = 8'h00;
    mem[974] = 8'h00;
    mem[975] = 8'h00;
    mem[976] = 8'h00;
    mem[977] = 8'h00;
    mem[978] = 8'h00;
    mem[979] = 8'h00;
    mem[980] = 8'h00;
    mem[981] = 8'h00;
    mem[982] = 8'h00;
    mem[983] = 8'h00;
    mem[984] = 8'h00;
    mem[985] = 8'h00;
    mem[986] = 8'h00;
    mem[987] = 8'h00;
    mem[988] = 8'h00;
    mem[989] = 8'h00;
    mem[990] = 8'h00;
    mem[991] = 8'h00;
    mem[992] = 8'h00;
    mem[993] = 8'h00;
    mem[994] = 8'h00;
    mem[995] = 8'h00;
    mem[996] = 8'h00;
    mem[997] = 8'h00;
    mem[998] = 8'h00;
    mem[999] = 8'h00;
    mem[1000] = 8'h00;
    mem[1001] = 8'h00;
    mem[1002] = 8'h00;
    mem[1003] = 8'h00;
    mem[1004] = 8'h00;
    mem[1005] = 8'h00;
    mem[1006] = 8'h00;
    mem[1007] = 8'h00;
    mem[1008] = 8'h00;
    mem[1009] = 8'h00;
    mem[1010] = 8'h00;
    mem[1011] = 8'h00;
    mem[1012] = 8'h00;
    mem[1013] = 8'h00;
    mem[1014] = 8'h00;
    mem[1015] = 8'h00;
    mem[1016] = 8'h00;
    mem[1017] = 8'h00;
    mem[1018] = 8'h00;
    mem[1019] = 8'h00;
    mem[1020] = 8'h00;
    mem[1021] = 8'h00;
    mem[1022] = 8'h00;
    mem[1023] = 8'h00;
    mem[1024] = 8'h00;
    mem[1025] = 8'h00;
    mem[1026] = 8'h00;
    mem[1027] = 8'h00;
    mem[1028] = 8'h00;
    mem[1029] = 8'h00;
    mem[1030] = 8'h00;
    mem[1031] = 8'h00;
    mem[1032] = 8'h00;
    mem[1033] = 8'h00;
    mem[1034] = 8'h00;
    mem[1035] = 8'h00;
    mem[1036] = 8'h00;
    mem[1037] = 8'h00;
    mem[1038] = 8'h00;
    mem[1039] = 8'h00;
    mem[1040] = 8'h00;
    mem[1041] = 8'h00;
    mem[1042] = 8'h00;
    mem[1043] = 8'h00;
    mem[1044] = 8'h00;
    mem[1045] = 8'h00;
    mem[1046] = 8'h00;
    mem[1047] = 8'h00;
    mem[1048] = 8'h00;
    mem[1049] = 8'h00;
    mem[1050] = 8'h00;
    mem[1051] = 8'h00;
    mem[1052] = 8'h00;
    mem[1053] = 8'h00;
    mem[1054] = 8'h00;
    mem[1055] = 8'h00;
    mem[1056] = 8'h00;
    mem[1057] = 8'h00;
    mem[1058] = 8'h00;
    mem[1059] = 8'h00;
    mem[1060] = 8'h00;
    mem[1061] = 8'h00;
    mem[1062] = 8'h00;
    mem[1063] = 8'h00;
    mem[1064] = 8'h00;
    mem[1065] = 8'h00;
    mem[1066] = 8'h00;
    mem[1067] = 8'h00;
    mem[1068] = 8'h00;
    mem[1069] = 8'h00;
    mem[1070] = 8'h00;
    mem[1071] = 8'h00;
    mem[1072] = 8'h00;
    mem[1073] = 8'h00;
    mem[1074] = 8'h80;
    mem[1075] = 8'hff;
    mem[1076] = 8'h02;
    mem[1077] = 8'h00;
    mem[1078] = 8'h00;
    mem[1079] = 8'h00;
    mem[1080] = 8'h00;
    mem[1081] = 8'h00;
    mem[1082] = 8'h00;
    mem[1083] = 8'h00;
    mem[1084] = 8'h00;
    mem[1085] = 8'h00;
    mem[1086] = 8'h00;
    mem[1087] = 8'h00;
    mem[1088] = 8'h00;
    mem[1089] = 8'h00;
    mem[1090] = 8'hff;
    mem[1091] = 8'hff;
    mem[1092] = 8'hff;
    mem[1093] = 8'h01;
    mem[1094] = 8'h00;
    mem[1095] = 8'h00;
    mem[1096] = 8'h00;
    mem[1097] = 8'hf8;
    mem[1098] = 8'hff;
    mem[1099] = 8'hff;
    mem[1100] = 8'h07;
    mem[1101] = 8'h00;
    mem[1102] = 8'h00;
    mem[1103] = 8'h00;
    mem[1104] = 8'h00;
    mem[1105] = 8'hc0;
    mem[1106] = 8'hff;
    mem[1107] = 8'hff;
    mem[1108] = 8'hff;
    mem[1109] = 8'h0f;
    mem[1110] = 8'h00;
    mem[1111] = 8'h00;
    mem[1112] = 8'h00;
    mem[1113] = 8'hfe;
    mem[1114] = 8'hff;
    mem[1115] = 8'hff;
    mem[1116] = 8'h7f;
    mem[1117] = 8'h00;
    mem[1118] = 8'h00;
    mem[1119] = 8'h00;
    mem[1120] = 8'h00;
    mem[1121] = 8'he0;
    mem[1122] = 8'hff;
    mem[1123] = 8'hff;
    mem[1124] = 8'hff;
    mem[1125] = 8'h3f;
    mem[1126] = 8'h00;
    mem[1127] = 8'h00;
    mem[1128] = 8'h00;
    mem[1129] = 8'hff;
    mem[1130] = 8'hff;
    mem[1131] = 8'hff;
    mem[1132] = 8'hff;
    mem[1133] = 8'h01;
    mem[1134] = 8'h00;
    mem[1135] = 8'h00;
    mem[1136] = 8'h00;
    mem[1137] = 8'he0;
    mem[1138] = 8'hff;
    mem[1139] = 8'hff;
    mem[1140] = 8'hff;
    mem[1141] = 8'hff;
    mem[1142] = 8'h00;
    mem[1143] = 8'h00;
    mem[1144] = 8'h80;
    mem[1145] = 8'hff;
    mem[1146] = 8'hff;
    mem[1147] = 8'hff;
    mem[1148] = 8'hff;
    mem[1149] = 8'h07;
    mem[1150] = 8'h00;
    mem[1151] = 8'h00;
    mem[1152] = 8'h00;
    mem[1153] = 8'hf0;
    mem[1154] = 8'hff;
    mem[1155] = 8'hff;
    mem[1156] = 8'hff;
    mem[1157] = 8'hff;
    mem[1158] = 8'h03;
    mem[1159] = 8'h00;
    mem[1160] = 8'h80;
    mem[1161] = 8'hff;
    mem[1162] = 8'hff;
    mem[1163] = 8'hff;
    mem[1164] = 8'hff;
    mem[1165] = 8'h1f;
    mem[1166] = 8'h00;
    mem[1167] = 8'h00;
    mem[1168] = 8'h00;
    mem[1169] = 8'hf0;
    mem[1170] = 8'hff;
    mem[1171] = 8'hff;
    mem[1172] = 8'hff;
    mem[1173] = 8'hff;
    mem[1174] = 8'h07;
    mem[1175] = 8'h00;
    mem[1176] = 8'h80;
    mem[1177] = 8'hff;
    mem[1178] = 8'hff;
    mem[1179] = 8'hff;
    mem[1180] = 8'hff;
    mem[1181] = 8'h3f;
    mem[1182] = 8'h00;
    mem[1183] = 8'h00;
    mem[1184] = 8'h00;
    mem[1185] = 8'hf0;
    mem[1186] = 8'hff;
    mem[1187] = 8'hff;
    mem[1188] = 8'hff;
    mem[1189] = 8'hff;
    mem[1190] = 8'h0f;
    mem[1191] = 8'h00;
    mem[1192] = 8'hc0;
    mem[1193] = 8'hff;
    mem[1194] = 8'hff;
    mem[1195] = 8'hff;
    mem[1196] = 8'hff;
    mem[1197] = 8'h7f;
    mem[1198] = 8'h00;
    mem[1199] = 8'h00;
    mem[1200] = 8'h00;
    mem[1201] = 8'hf0;
    mem[1202] = 8'hff;
    mem[1203] = 8'hff;
    mem[1204] = 8'hff;
    mem[1205] = 8'hff;
    mem[1206] = 8'h1f;
    mem[1207] = 8'h00;
    mem[1208] = 8'hc0;
    mem[1209] = 8'hff;
    mem[1210] = 8'hff;
    mem[1211] = 8'hff;
    mem[1212] = 8'hff;
    mem[1213] = 8'hff;
    mem[1214] = 8'h00;
    mem[1215] = 8'h00;
    mem[1216] = 8'h00;
    mem[1217] = 8'hf0;
    mem[1218] = 8'hff;
    mem[1219] = 8'hff;
    mem[1220] = 8'hff;
    mem[1221] = 8'hff;
    mem[1222] = 8'h3f;
    mem[1223] = 8'h00;
    mem[1224] = 8'hc0;
    mem[1225] = 8'hff;
    mem[1226] = 8'hff;
    mem[1227] = 8'hff;
    mem[1228] = 8'hff;
    mem[1229] = 8'hff;
    mem[1230] = 8'h01;
    mem[1231] = 8'h00;
    mem[1232] = 8'h00;
    mem[1233] = 8'hf0;
    mem[1234] = 8'hff;
    mem[1235] = 8'hff;
    mem[1236] = 8'hff;
    mem[1237] = 8'hff;
    mem[1238] = 8'h7f;
    mem[1239] = 8'h00;
    mem[1240] = 8'hc0;
    mem[1241] = 8'hff;
    mem[1242] = 8'hff;
    mem[1243] = 8'hff;
    mem[1244] = 8'hff;
    mem[1245] = 8'hff;
    mem[1246] = 8'h03;
    mem[1247] = 8'h00;
    mem[1248] = 8'h00;
    mem[1249] = 8'hf0;
    mem[1250] = 8'hff;
    mem[1251] = 8'hff;
    mem[1252] = 8'hff;
    mem[1253] = 8'hff;
    mem[1254] = 8'hff;
    mem[1255] = 8'h00;
    mem[1256] = 8'hc0;
    mem[1257] = 8'hff;
    mem[1258] = 8'hff;
    mem[1259] = 8'hff;
    mem[1260] = 8'hff;
    mem[1261] = 8'hff;
    mem[1262] = 8'h07;
    mem[1263] = 8'h00;
    mem[1264] = 8'h00;
    mem[1265] = 8'hf0;
    mem[1266] = 8'hff;
    mem[1267] = 8'hff;
    mem[1268] = 8'hff;
    mem[1269] = 8'hff;
    mem[1270] = 8'hff;
    mem[1271] = 8'h00;
    mem[1272] = 8'hc0;
    mem[1273] = 8'hff;
    mem[1274] = 8'hff;
    mem[1275] = 8'hff;
    mem[1276] = 8'hff;
    mem[1277] = 8'hff;
    mem[1278] = 8'h07;
    mem[1279] = 8'h00;
    mem[1280] = 8'h00;
    mem[1281] = 8'hf0;
    mem[1282] = 8'hff;
    mem[1283] = 8'hff;
    mem[1284] = 8'hff;
    mem[1285] = 8'hff;
    mem[1286] = 8'hff;
    mem[1287] = 8'h01;
    mem[1288] = 8'hc0;
    mem[1289] = 8'hff;
    mem[1290] = 8'hff;
    mem[1291] = 8'hff;
    mem[1292] = 8'hff;
    mem[1293] = 8'hff;
    mem[1294] = 8'h0f;
    mem[1295] = 8'h00;
    mem[1296] = 8'h00;
    mem[1297] = 8'hf0;
    mem[1298] = 8'hff;
    mem[1299] = 8'hff;
    mem[1300] = 8'hff;
    mem[1301] = 8'hff;
    mem[1302] = 8'hff;
    mem[1303] = 8'h01;
    mem[1304] = 8'hc0;
    mem[1305] = 8'hff;
    mem[1306] = 8'hff;
    mem[1307] = 8'hff;
    mem[1308] = 8'hff;
    mem[1309] = 8'hff;
    mem[1310] = 8'h0f;
    mem[1311] = 8'h00;
    mem[1312] = 8'h00;
    mem[1313] = 8'hf0;
    mem[1314] = 8'hff;
    mem[1315] = 8'hff;
    mem[1316] = 8'hff;
    mem[1317] = 8'hff;
    mem[1318] = 8'hff;
    mem[1319] = 8'h03;
    mem[1320] = 8'hc0;
    mem[1321] = 8'hff;
    mem[1322] = 8'hff;
    mem[1323] = 8'hff;
    mem[1324] = 8'hff;
    mem[1325] = 8'hff;
    mem[1326] = 8'h1f;
    mem[1327] = 8'h00;
    mem[1328] = 8'h00;
    mem[1329] = 8'hf0;
    mem[1330] = 8'hff;
    mem[1331] = 8'hff;
    mem[1332] = 8'hff;
    mem[1333] = 8'hff;
    mem[1334] = 8'hff;
    mem[1335] = 8'h03;
    mem[1336] = 8'hc0;
    mem[1337] = 8'hff;
    mem[1338] = 8'hff;
    mem[1339] = 8'hff;
    mem[1340] = 8'hff;
    mem[1341] = 8'hff;
    mem[1342] = 8'h1f;
    mem[1343] = 8'h00;
    mem[1344] = 8'h00;
    mem[1345] = 8'hf0;
    mem[1346] = 8'hff;
    mem[1347] = 8'hff;
    mem[1348] = 8'hff;
    mem[1349] = 8'hff;
    mem[1350] = 8'hff;
    mem[1351] = 8'h07;
    mem[1352] = 8'hc0;
    mem[1353] = 8'hff;
    mem[1354] = 8'hff;
    mem[1355] = 8'hff;
    mem[1356] = 8'hff;
    mem[1357] = 8'hff;
    mem[1358] = 8'h3f;
    mem[1359] = 8'h00;
    mem[1360] = 8'h00;
    mem[1361] = 8'hf0;
    mem[1362] = 8'hff;
    mem[1363] = 8'hff;
    mem[1364] = 8'hff;
    mem[1365] = 8'hff;
    mem[1366] = 8'hff;
    mem[1367] = 8'h07;
    mem[1368] = 8'hc0;
    mem[1369] = 8'hff;
    mem[1370] = 8'hff;
    mem[1371] = 8'hff;
    mem[1372] = 8'hff;
    mem[1373] = 8'hff;
    mem[1374] = 8'h3f;
    mem[1375] = 8'h00;
    mem[1376] = 8'h00;
    mem[1377] = 8'hf0;
    mem[1378] = 8'hff;
    mem[1379] = 8'hff;
    mem[1380] = 8'hff;
    mem[1381] = 8'hff;
    mem[1382] = 8'hff;
    mem[1383] = 8'h07;
    mem[1384] = 8'hc0;
    mem[1385] = 8'hff;
    mem[1386] = 8'hff;
    mem[1387] = 8'hff;
    mem[1388] = 8'hff;
    mem[1389] = 8'hff;
    mem[1390] = 8'h3f;
    mem[1391] = 8'h00;
    mem[1392] = 8'h00;
    mem[1393] = 8'hf0;
    mem[1394] = 8'hff;
    mem[1395] = 8'hff;
    mem[1396] = 8'hff;
    mem[1397] = 8'hff;
    mem[1398] = 8'hff;
    mem[1399] = 8'h0f;
    mem[1400] = 8'hc0;
    mem[1401] = 8'hff;
    mem[1402] = 8'hff;
    mem[1403] = 8'hff;
    mem[1404] = 8'hff;
    mem[1405] = 8'hff;
    mem[1406] = 8'h3f;
    mem[1407] = 8'h00;
    mem[1408] = 8'h00;
    mem[1409] = 8'hf0;
    mem[1410] = 8'hff;
    mem[1411] = 8'hff;
    mem[1412] = 8'hff;
    mem[1413] = 8'hff;
    mem[1414] = 8'hff;
    mem[1415] = 8'h0f;
    mem[1416] = 8'hc0;
    mem[1417] = 8'hff;
    mem[1418] = 8'hff;
    mem[1419] = 8'hff;
    mem[1420] = 8'hff;
    mem[1421] = 8'hff;
    mem[1422] = 8'h7f;
    mem[1423] = 8'h00;
    mem[1424] = 8'h00;
    mem[1425] = 8'hf0;
    mem[1426] = 8'hff;
    mem[1427] = 8'hff;
    mem[1428] = 8'hff;
    mem[1429] = 8'hff;
    mem[1430] = 8'hff;
    mem[1431] = 8'h0f;
    mem[1432] = 8'hc0;
    mem[1433] = 8'hff;
    mem[1434] = 8'hff;
    mem[1435] = 8'hff;
    mem[1436] = 8'hff;
    mem[1437] = 8'hff;
    mem[1438] = 8'h7f;
    mem[1439] = 8'h00;
    mem[1440] = 8'h00;
    mem[1441] = 8'hf0;
    mem[1442] = 8'hff;
    mem[1443] = 8'hff;
    mem[1444] = 8'hff;
    mem[1445] = 8'hff;
    mem[1446] = 8'hff;
    mem[1447] = 8'h0f;
    mem[1448] = 8'hc0;
    mem[1449] = 8'hff;
    mem[1450] = 8'hff;
    mem[1451] = 8'hff;
    mem[1452] = 8'hff;
    mem[1453] = 8'hff;
    mem[1454] = 8'h7f;
    mem[1455] = 8'h00;
    mem[1456] = 8'h00;
    mem[1457] = 8'hf0;
    mem[1458] = 8'hff;
    mem[1459] = 8'hff;
    mem[1460] = 8'hff;
    mem[1461] = 8'hff;
    mem[1462] = 8'hff;
    mem[1463] = 8'h0f;
    mem[1464] = 8'hc0;
    mem[1465] = 8'hff;
    mem[1466] = 8'hff;
    mem[1467] = 8'hff;
    mem[1468] = 8'hff;
    mem[1469] = 8'hff;
    mem[1470] = 8'h7f;
    mem[1471] = 8'h00;
    mem[1472] = 8'h00;
    mem[1473] = 8'hf0;
    mem[1474] = 8'hff;
    mem[1475] = 8'hff;
    mem[1476] = 8'hff;
    mem[1477] = 8'hff;
    mem[1478] = 8'hff;
    mem[1479] = 8'h0f;
    mem[1480] = 8'hc0;
    mem[1481] = 8'hff;
    mem[1482] = 8'hff;
    mem[1483] = 8'hff;
    mem[1484] = 8'hff;
    mem[1485] = 8'hff;
    mem[1486] = 8'h7f;
    mem[1487] = 8'h00;
    mem[1488] = 8'h00;
    mem[1489] = 8'hf0;
    mem[1490] = 8'hff;
    mem[1491] = 8'hff;
    mem[1492] = 8'hff;
    mem[1493] = 8'hff;
    mem[1494] = 8'hff;
    mem[1495] = 8'h0f;
    mem[1496] = 8'hc0;
    mem[1497] = 8'hff;
    mem[1498] = 8'hff;
    mem[1499] = 8'hff;
    mem[1500] = 8'hff;
    mem[1501] = 8'hff;
    mem[1502] = 8'h7f;
    mem[1503] = 8'h00;
    mem[1504] = 8'h00;
    mem[1505] = 8'hf0;
    mem[1506] = 8'hff;
    mem[1507] = 8'hff;
    mem[1508] = 8'hff;
    mem[1509] = 8'hff;
    mem[1510] = 8'hff;
    mem[1511] = 8'h0f;
    mem[1512] = 8'hc0;
    mem[1513] = 8'hff;
    mem[1514] = 8'hff;
    mem[1515] = 8'hff;
    mem[1516] = 8'hff;
    mem[1517] = 8'hff;
    mem[1518] = 8'h7f;
    mem[1519] = 8'h00;
    mem[1520] = 8'h00;
    mem[1521] = 8'hf0;
    mem[1522] = 8'hff;
    mem[1523] = 8'hff;
    mem[1524] = 8'hff;
    mem[1525] = 8'hff;
    mem[1526] = 8'hff;
    mem[1527] = 8'h0f;
    mem[1528] = 8'hc0;
    mem[1529] = 8'hff;
    mem[1530] = 8'hff;
    mem[1531] = 8'hff;
    mem[1532] = 8'hff;
    mem[1533] = 8'hff;
    mem[1534] = 8'h7f;
    mem[1535] = 8'h00;
    mem[1536] = 8'h00;
    mem[1537] = 8'hf0;
    mem[1538] = 8'hff;
    mem[1539] = 8'hff;
    mem[1540] = 8'hff;
    mem[1541] = 8'hff;
    mem[1542] = 8'hff;
    mem[1543] = 8'h0f;
    mem[1544] = 8'hc0;
    mem[1545] = 8'hff;
    mem[1546] = 8'hff;
    mem[1547] = 8'hff;
    mem[1548] = 8'hff;
    mem[1549] = 8'hff;
    mem[1550] = 8'h7f;
    mem[1551] = 8'h00;
    mem[1552] = 8'h00;
    mem[1553] = 8'hf0;
    mem[1554] = 8'hff;
    mem[1555] = 8'hff;
    mem[1556] = 8'hff;
    mem[1557] = 8'hff;
    mem[1558] = 8'hff;
    mem[1559] = 8'h0f;
    mem[1560] = 8'hc0;
    mem[1561] = 8'hff;
    mem[1562] = 8'hff;
    mem[1563] = 8'hff;
    mem[1564] = 8'hff;
    mem[1565] = 8'hff;
    mem[1566] = 8'h7f;
    mem[1567] = 8'h00;
    mem[1568] = 8'h00;
    mem[1569] = 8'hf0;
    mem[1570] = 8'hff;
    mem[1571] = 8'hff;
    mem[1572] = 8'hff;
    mem[1573] = 8'hff;
    mem[1574] = 8'hff;
    mem[1575] = 8'h0f;
    mem[1576] = 8'hc0;
    mem[1577] = 8'hff;
    mem[1578] = 8'hff;
    mem[1579] = 8'hff;
    mem[1580] = 8'hff;
    mem[1581] = 8'hff;
    mem[1582] = 8'h7f;
    mem[1583] = 8'h00;
    mem[1584] = 8'h00;
    mem[1585] = 8'hf0;
    mem[1586] = 8'hff;
    mem[1587] = 8'hff;
    mem[1588] = 8'hff;
    mem[1589] = 8'hff;
    mem[1590] = 8'hff;
    mem[1591] = 8'h0f;
    mem[1592] = 8'hc0;
    mem[1593] = 8'hff;
    mem[1594] = 8'hff;
    mem[1595] = 8'hff;
    mem[1596] = 8'hff;
    mem[1597] = 8'hff;
    mem[1598] = 8'h7f;
    mem[1599] = 8'h00;
    mem[1600] = 8'h00;
    mem[1601] = 8'hf0;
    mem[1602] = 8'hff;
    mem[1603] = 8'hff;
    mem[1604] = 8'hff;
    mem[1605] = 8'hff;
    mem[1606] = 8'hff;
    mem[1607] = 8'h0f;
    mem[1608] = 8'hc0;
    mem[1609] = 8'hff;
    mem[1610] = 8'hff;
    mem[1611] = 8'hff;
    mem[1612] = 8'hff;
    mem[1613] = 8'hff;
    mem[1614] = 8'h7f;
    mem[1615] = 8'h00;
    mem[1616] = 8'h00;
    mem[1617] = 8'hf0;
    mem[1618] = 8'hff;
    mem[1619] = 8'hff;
    mem[1620] = 8'hff;
    mem[1621] = 8'hff;
    mem[1622] = 8'hff;
    mem[1623] = 8'h07;
    mem[1624] = 8'hc0;
    mem[1625] = 8'hff;
    mem[1626] = 8'hff;
    mem[1627] = 8'hff;
    mem[1628] = 8'hff;
    mem[1629] = 8'hff;
    mem[1630] = 8'h3f;
    mem[1631] = 8'h00;
    mem[1632] = 8'h00;
    mem[1633] = 8'hf0;
    mem[1634] = 8'hff;
    mem[1635] = 8'hff;
    mem[1636] = 8'hff;
    mem[1637] = 8'hff;
    mem[1638] = 8'hff;
    mem[1639] = 8'h07;
    mem[1640] = 8'hc0;
    mem[1641] = 8'hff;
    mem[1642] = 8'hff;
    mem[1643] = 8'hff;
    mem[1644] = 8'hff;
    mem[1645] = 8'hff;
    mem[1646] = 8'h3f;
    mem[1647] = 8'h00;
    mem[1648] = 8'h00;
    mem[1649] = 8'hf0;
    mem[1650] = 8'hff;
    mem[1651] = 8'hff;
    mem[1652] = 8'hff;
    mem[1653] = 8'hff;
    mem[1654] = 8'hff;
    mem[1655] = 8'h07;
    mem[1656] = 8'hc0;
    mem[1657] = 8'hff;
    mem[1658] = 8'hff;
    mem[1659] = 8'hff;
    mem[1660] = 8'hff;
    mem[1661] = 8'hff;
    mem[1662] = 8'h3f;
    mem[1663] = 8'h00;
    mem[1664] = 8'h00;
    mem[1665] = 8'hf0;
    mem[1666] = 8'hff;
    mem[1667] = 8'hff;
    mem[1668] = 8'hff;
    mem[1669] = 8'hff;
    mem[1670] = 8'hff;
    mem[1671] = 8'h07;
    mem[1672] = 8'hc0;
    mem[1673] = 8'hff;
    mem[1674] = 8'hff;
    mem[1675] = 8'hff;
    mem[1676] = 8'hff;
    mem[1677] = 8'hff;
    mem[1678] = 8'h3f;
    mem[1679] = 8'h00;
    mem[1680] = 8'h00;
    mem[1681] = 8'hf0;
    mem[1682] = 8'hff;
    mem[1683] = 8'hff;
    mem[1684] = 8'hff;
    mem[1685] = 8'hff;
    mem[1686] = 8'hff;
    mem[1687] = 8'h03;
    mem[1688] = 8'hc0;
    mem[1689] = 8'hff;
    mem[1690] = 8'hff;
    mem[1691] = 8'hff;
    mem[1692] = 8'hff;
    mem[1693] = 8'hff;
    mem[1694] = 8'h1f;
    mem[1695] = 8'h00;
    mem[1696] = 8'h00;
    mem[1697] = 8'hf0;
    mem[1698] = 8'hff;
    mem[1699] = 8'hff;
    mem[1700] = 8'hff;
    mem[1701] = 8'hff;
    mem[1702] = 8'hff;
    mem[1703] = 8'h03;
    mem[1704] = 8'hc0;
    mem[1705] = 8'hff;
    mem[1706] = 8'hff;
    mem[1707] = 8'hff;
    mem[1708] = 8'hff;
    mem[1709] = 8'hff;
    mem[1710] = 8'h1f;
    mem[1711] = 8'h00;
    mem[1712] = 8'h00;
    mem[1713] = 8'hf0;
    mem[1714] = 8'hff;
    mem[1715] = 8'hff;
    mem[1716] = 8'hff;
    mem[1717] = 8'hff;
    mem[1718] = 8'hff;
    mem[1719] = 8'h01;
    mem[1720] = 8'hc0;
    mem[1721] = 8'hff;
    mem[1722] = 8'hff;
    mem[1723] = 8'hff;
    mem[1724] = 8'hff;
    mem[1725] = 8'hff;
    mem[1726] = 8'h0f;
    mem[1727] = 8'h00;
    mem[1728] = 8'h00;
    mem[1729] = 8'hf0;
    mem[1730] = 8'hff;
    mem[1731] = 8'hff;
    mem[1732] = 8'hff;
    mem[1733] = 8'hff;
    mem[1734] = 8'hff;
    mem[1735] = 8'h01;
    mem[1736] = 8'hc0;
    mem[1737] = 8'hff;
    mem[1738] = 8'hff;
    mem[1739] = 8'hff;
    mem[1740] = 8'hff;
    mem[1741] = 8'hff;
    mem[1742] = 8'h0f;
    mem[1743] = 8'h00;
    mem[1744] = 8'h00;
    mem[1745] = 8'hf0;
    mem[1746] = 8'hff;
    mem[1747] = 8'hff;
    mem[1748] = 8'hff;
    mem[1749] = 8'hff;
    mem[1750] = 8'hff;
    mem[1751] = 8'h00;
    mem[1752] = 8'hc0;
    mem[1753] = 8'hff;
    mem[1754] = 8'hff;
    mem[1755] = 8'hff;
    mem[1756] = 8'hff;
    mem[1757] = 8'hff;
    mem[1758] = 8'h07;
    mem[1759] = 8'h00;
    mem[1760] = 8'h00;
    mem[1761] = 8'hf0;
    mem[1762] = 8'hff;
    mem[1763] = 8'hff;
    mem[1764] = 8'hff;
    mem[1765] = 8'hff;
    mem[1766] = 8'h7f;
    mem[1767] = 8'h00;
    mem[1768] = 8'hc0;
    mem[1769] = 8'hff;
    mem[1770] = 8'hff;
    mem[1771] = 8'hff;
    mem[1772] = 8'hff;
    mem[1773] = 8'hff;
    mem[1774] = 8'h03;
    mem[1775] = 8'h00;
    mem[1776] = 8'h00;
    mem[1777] = 8'hf0;
    mem[1778] = 8'hff;
    mem[1779] = 8'hff;
    mem[1780] = 8'hff;
    mem[1781] = 8'hff;
    mem[1782] = 8'h7f;
    mem[1783] = 8'h00;
    mem[1784] = 8'hc0;
    mem[1785] = 8'hff;
    mem[1786] = 8'hff;
    mem[1787] = 8'hff;
    mem[1788] = 8'hff;
    mem[1789] = 8'hff;
    mem[1790] = 8'h01;
    mem[1791] = 8'h00;
    mem[1792] = 8'h00;
    mem[1793] = 8'hf0;
    mem[1794] = 8'hff;
    mem[1795] = 8'hff;
    mem[1796] = 8'hff;
    mem[1797] = 8'hff;
    mem[1798] = 8'h3f;
    mem[1799] = 8'h00;
    mem[1800] = 8'hc0;
    mem[1801] = 8'hff;
    mem[1802] = 8'hff;
    mem[1803] = 8'hff;
    mem[1804] = 8'hff;
    mem[1805] = 8'hff;
    mem[1806] = 8'h01;
    mem[1807] = 8'h00;
    mem[1808] = 8'h00;
    mem[1809] = 8'hf0;
    mem[1810] = 8'hff;
    mem[1811] = 8'hff;
    mem[1812] = 8'hff;
    mem[1813] = 8'hff;
    mem[1814] = 8'h1f;
    mem[1815] = 8'h00;
    mem[1816] = 8'hc0;
    mem[1817] = 8'hff;
    mem[1818] = 8'hff;
    mem[1819] = 8'hff;
    mem[1820] = 8'hff;
    mem[1821] = 8'hff;
    mem[1822] = 8'h00;
    mem[1823] = 8'h00;
    mem[1824] = 8'h00;
    mem[1825] = 8'hf0;
    mem[1826] = 8'hff;
    mem[1827] = 8'hff;
    mem[1828] = 8'hff;
    mem[1829] = 8'hff;
    mem[1830] = 8'h0f;
    mem[1831] = 8'h00;
    mem[1832] = 8'h80;
    mem[1833] = 8'hff;
    mem[1834] = 8'hff;
    mem[1835] = 8'hff;
    mem[1836] = 8'hff;
    mem[1837] = 8'h7f;
    mem[1838] = 8'h00;
    mem[1839] = 8'h00;
    mem[1840] = 8'h00;
    mem[1841] = 8'hf0;
    mem[1842] = 8'hff;
    mem[1843] = 8'hff;
    mem[1844] = 8'hff;
    mem[1845] = 8'hff;
    mem[1846] = 8'h03;
    mem[1847] = 8'h00;
    mem[1848] = 8'h80;
    mem[1849] = 8'hff;
    mem[1850] = 8'hff;
    mem[1851] = 8'hff;
    mem[1852] = 8'hff;
    mem[1853] = 8'h1f;
    mem[1854] = 8'h00;
    mem[1855] = 8'h00;
    mem[1856] = 8'h00;
    mem[1857] = 8'hf0;
    mem[1858] = 8'hff;
    mem[1859] = 8'hff;
    mem[1860] = 8'hff;
    mem[1861] = 8'hff;
    mem[1862] = 8'h01;
    mem[1863] = 8'h00;
    mem[1864] = 8'h80;
    mem[1865] = 8'hff;
    mem[1866] = 8'hff;
    mem[1867] = 8'hff;
    mem[1868] = 8'hff;
    mem[1869] = 8'h0f;
    mem[1870] = 8'h00;
    mem[1871] = 8'h00;
    mem[1872] = 8'h00;
    mem[1873] = 8'he0;
    mem[1874] = 8'hff;
    mem[1875] = 8'hff;
    mem[1876] = 8'hff;
    mem[1877] = 8'hff;
    mem[1878] = 8'h00;
    mem[1879] = 8'h00;
    mem[1880] = 8'h00;
    mem[1881] = 8'hff;
    mem[1882] = 8'hff;
    mem[1883] = 8'hff;
    mem[1884] = 8'hff;
    mem[1885] = 8'h07;
    mem[1886] = 8'h00;
    mem[1887] = 8'h00;
    mem[1888] = 8'h00;
    mem[1889] = 8'hc0;
    mem[1890] = 8'hff;
    mem[1891] = 8'hff;
    mem[1892] = 8'hff;
    mem[1893] = 8'h3f;
    mem[1894] = 8'h00;
    mem[1895] = 8'h00;
    mem[1896] = 8'h00;
    mem[1897] = 8'hfe;
    mem[1898] = 8'hff;
    mem[1899] = 8'hff;
    mem[1900] = 8'hff;
    mem[1901] = 8'h01;
    mem[1902] = 8'h00;
    mem[1903] = 8'h00;
    mem[1904] = 8'h00;
    mem[1905] = 8'h80;
    mem[1906] = 8'hff;
    mem[1907] = 8'hff;
    mem[1908] = 8'hff;
    mem[1909] = 8'h07;
    mem[1910] = 8'h00;
    mem[1911] = 8'h00;
    mem[1912] = 8'h00;
    mem[1913] = 8'hfc;
    mem[1914] = 8'hff;
    mem[1915] = 8'hff;
    mem[1916] = 8'h3f;
    mem[1917] = 8'h00;
    mem[1918] = 8'h00;
    mem[1919] = 8'h00;
    mem[1920] = 8'h00;
    mem[1921] = 8'h00;
    mem[1922] = 8'hff;
    mem[1923] = 8'hff;
    mem[1924] = 8'hff;
    mem[1925] = 8'h00;
    mem[1926] = 8'h00;
    mem[1927] = 8'h00;
    mem[1928] = 8'h00;
    mem[1929] = 8'hf8;
    mem[1930] = 8'hff;
    mem[1931] = 8'hff;
    mem[1932] = 8'h03;
    mem[1933] = 8'h00;
    mem[1934] = 8'h00;
    mem[1935] = 8'h00;
    mem[1936] = 8'h00;
    mem[1937] = 8'h00;
    mem[1938] = 8'h00;
    mem[1939] = 8'h00;
    mem[1940] = 8'h00;
    mem[1941] = 8'h00;
    mem[1942] = 8'h00;
    mem[1943] = 8'h00;
    mem[1944] = 8'h00;
    mem[1945] = 8'h00;
    mem[1946] = 8'h00;
    mem[1947] = 8'h00;
    mem[1948] = 8'h00;
    mem[1949] = 8'h00;
    mem[1950] = 8'h00;
    mem[1951] = 8'h00;
    mem[1952] = 8'h00;
    mem[1953] = 8'h00;
    mem[1954] = 8'h00;
    mem[1955] = 8'h00;
    mem[1956] = 8'h00;
    mem[1957] = 8'h00;
    mem[1958] = 8'h00;
    mem[1959] = 8'h00;
    mem[1960] = 8'h00;
    mem[1961] = 8'h00;
    mem[1962] = 8'h00;
    mem[1963] = 8'h00;
    mem[1964] = 8'h00;
    mem[1965] = 8'h00;
    mem[1966] = 8'h00;
    mem[1967] = 8'h00;
    mem[1968] = 8'h00;
    mem[1969] = 8'h00;
    mem[1970] = 8'h00;
    mem[1971] = 8'h00;
    mem[1972] = 8'h00;
    mem[1973] = 8'h00;
    mem[1974] = 8'h00;
    mem[1975] = 8'h00;
    mem[1976] = 8'h00;
    mem[1977] = 8'h00;
    mem[1978] = 8'h00;
    mem[1979] = 8'h00;
    mem[1980] = 8'h00;
    mem[1981] = 8'h00;
    mem[1982] = 8'h00;
    mem[1983] = 8'h00;
    mem[1984] = 8'h00;
    mem[1985] = 8'h00;
    mem[1986] = 8'h00;
    mem[1987] = 8'h00;
    mem[1988] = 8'h00;
    mem[1989] = 8'h00;
    mem[1990] = 8'h00;
    mem[1991] = 8'h00;
    mem[1992] = 8'h00;
    mem[1993] = 8'h00;
    mem[1994] = 8'h00;
    mem[1995] = 8'h00;
    mem[1996] = 8'h00;
    mem[1997] = 8'h00;
    mem[1998] = 8'h00;
    mem[1999] = 8'h00;
    mem[2000] = 8'h00;
    mem[2001] = 8'h00;
    mem[2002] = 8'h00;
    mem[2003] = 8'h00;
    mem[2004] = 8'h00;
    mem[2005] = 8'h00;
    mem[2006] = 8'h00;
    mem[2007] = 8'h00;
    mem[2008] = 8'h00;
    mem[2009] = 8'h00;
    mem[2010] = 8'h00;
    mem[2011] = 8'h00;
    mem[2012] = 8'h00;
    mem[2013] = 8'h00;
    mem[2014] = 8'h00;
    mem[2015] = 8'h00;
    mem[2016] = 8'h00;
    mem[2017] = 8'h00;
    mem[2018] = 8'h00;
    mem[2019] = 8'h00;
    mem[2020] = 8'h00;
    mem[2021] = 8'h00;
    mem[2022] = 8'h00;
    mem[2023] = 8'h00;
    mem[2024] = 8'h00;
    mem[2025] = 8'h00;
    mem[2026] = 8'h00;
    mem[2027] = 8'h00;
    mem[2028] = 8'h00;
    mem[2029] = 8'h00;
    mem[2030] = 8'h00;
    mem[2031] = 8'h00;
    mem[2032] = 8'h00;
    mem[2033] = 8'h00;
    mem[2034] = 8'h00;
    mem[2035] = 8'h00;
    mem[2036] = 8'h00;
    mem[2037] = 8'h00;
    mem[2038] = 8'h00;
    mem[2039] = 8'h00;
    mem[2040] = 8'h00;
    mem[2041] = 8'h00;
    mem[2042] = 8'h00;
    mem[2043] = 8'h00;
    mem[2044] = 8'h00;
    mem[2045] = 8'h00;
    mem[2046] = 8'h00;
    mem[2047] = 8'h00;
  end

  wire [10:0] addr = {y[6:0], x[6:3]};
  assign pixel = mem[addr][x&7];

endmodule
