//`timescale 1ns / 1ps
module bitmap_rom_sk (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire pixel
);

  reg [7:0] mem[2047:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'he0;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'hf0;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'hf0;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h7c;
    mem[50] = 8'h1e;
    mem[51] = 8'h7c;
    mem[52] = 8'h80;
    mem[53] = 8'h8f;
    mem[54] = 8'h7b;
    mem[55] = 8'he0;
    mem[56] = 8'h70;
    mem[57] = 8'hf0;
    mem[58] = 8'hf8;
    mem[59] = 8'h1c;
    mem[60] = 8'hc0;
    mem[61] = 8'h03;
    mem[62] = 8'h3e;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'hfe;
    mem[66] = 8'h1f;
    mem[67] = 8'hff;
    mem[68] = 8'hc0;
    mem[69] = 8'hdf;
    mem[70] = 8'hff;
    mem[71] = 8'hf0;
    mem[72] = 8'h78;
    mem[73] = 8'hf8;
    mem[74] = 8'hfc;
    mem[75] = 8'h3d;
    mem[76] = 8'hc0;
    mem[77] = 8'hc3;
    mem[78] = 8'hff;
    mem[79] = 8'h01;
    mem[80] = 8'h00;
    mem[81] = 8'h0f;
    mem[82] = 8'h1e;
    mem[83] = 8'he7;
    mem[84] = 8'he1;
    mem[85] = 8'hf9;
    mem[86] = 8'hf3;
    mem[87] = 8'he0;
    mem[88] = 8'h78;
    mem[89] = 8'hf0;
    mem[90] = 8'h1e;
    mem[91] = 8'h1c;
    mem[92] = 8'hc0;
    mem[93] = 8'hc3;
    mem[94] = 8'hc3;
    mem[95] = 8'h01;
    mem[96] = 8'h80;
    mem[97] = 8'h07;
    mem[98] = 8'h1e;
    mem[99] = 8'hc3;
    mem[100] = 8'he3;
    mem[101] = 8'he0;
    mem[102] = 8'hf3;
    mem[103] = 8'he0;
    mem[104] = 8'h78;
    mem[105] = 8'hf0;
    mem[106] = 8'h1e;
    mem[107] = 8'h1c;
    mem[108] = 8'hc0;
    mem[109] = 8'he1;
    mem[110] = 8'hc1;
    mem[111] = 8'h01;
    mem[112] = 8'h00;
    mem[113] = 8'h0f;
    mem[114] = 8'h1e;
    mem[115] = 8'h80;
    mem[116] = 8'he3;
    mem[117] = 8'hc0;
    mem[118] = 8'hf3;
    mem[119] = 8'he0;
    mem[120] = 8'h78;
    mem[121] = 8'hf0;
    mem[122] = 8'h1e;
    mem[123] = 8'h1c;
    mem[124] = 8'hc0;
    mem[125] = 8'he1;
    mem[126] = 8'hc1;
    mem[127] = 8'h01;
    mem[128] = 8'h00;
    mem[129] = 8'hfe;
    mem[130] = 8'h1e;
    mem[131] = 8'h80;
    mem[132] = 8'he7;
    mem[133] = 8'hc0;
    mem[134] = 8'hf3;
    mem[135] = 8'he0;
    mem[136] = 8'h78;
    mem[137] = 8'hf0;
    mem[138] = 8'hfc;
    mem[139] = 8'h1d;
    mem[140] = 8'hc0;
    mem[141] = 8'he1;
    mem[142] = 8'hc1;
    mem[143] = 8'h01;
    mem[144] = 8'h00;
    mem[145] = 8'hf8;
    mem[146] = 8'h1f;
    mem[147] = 8'h80;
    mem[148] = 8'he3;
    mem[149] = 8'hc0;
    mem[150] = 8'hf3;
    mem[151] = 8'he0;
    mem[152] = 8'hf8;
    mem[153] = 8'hf1;
    mem[154] = 8'hf0;
    mem[155] = 8'h1f;
    mem[156] = 8'hc0;
    mem[157] = 8'he1;
    mem[158] = 8'hc1;
    mem[159] = 8'h01;
    mem[160] = 8'h00;
    mem[161] = 8'h06;
    mem[162] = 8'h9e;
    mem[163] = 8'h81;
    mem[164] = 8'he3;
    mem[165] = 8'hc0;
    mem[166] = 8'he3;
    mem[167] = 8'he0;
    mem[168] = 8'hf8;
    mem[169] = 8'h79;
    mem[170] = 8'h0c;
    mem[171] = 8'h1c;
    mem[172] = 8'hc1;
    mem[173] = 8'he1;
    mem[174] = 8'hc1;
    mem[175] = 8'h01;
    mem[176] = 8'h00;
    mem[177] = 8'h0e;
    mem[178] = 8'hde;
    mem[179] = 8'hc1;
    mem[180] = 8'he3;
    mem[181] = 8'hc0;
    mem[182] = 8'hf3;
    mem[183] = 8'he0;
    mem[184] = 8'hf8;
    mem[185] = 8'h7f;
    mem[186] = 8'h1c;
    mem[187] = 8'h9c;
    mem[188] = 8'hc3;
    mem[189] = 8'he1;
    mem[190] = 8'hc1;
    mem[191] = 8'h01;
    mem[192] = 8'h00;
    mem[193] = 8'h9e;
    mem[194] = 8'hcf;
    mem[195] = 8'he7;
    mem[196] = 8'hf9;
    mem[197] = 8'hc0;
    mem[198] = 8'hf3;
    mem[199] = 8'hf0;
    mem[200] = 8'h7e;
    mem[201] = 8'h7e;
    mem[202] = 8'h3c;
    mem[203] = 8'h9e;
    mem[204] = 8'he7;
    mem[205] = 8'hf9;
    mem[206] = 8'hc1;
    mem[207] = 8'h03;
    mem[208] = 8'h00;
    mem[209] = 8'hf8;
    mem[210] = 8'h1f;
    mem[211] = 8'hff;
    mem[212] = 8'h70;
    mem[213] = 8'he0;
    mem[214] = 8'he3;
    mem[215] = 8'h3f;
    mem[216] = 8'h38;
    mem[217] = 8'hfe;
    mem[218] = 8'hf1;
    mem[219] = 8'h07;
    mem[220] = 8'hff;
    mem[221] = 8'he0;
    mem[222] = 8'he0;
    mem[223] = 8'h07;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h1c;
    mem[227] = 8'h00;
    mem[228] = 8'h00;
    mem[229] = 8'h00;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h00;
    mem[235] = 8'h00;
    mem[236] = 8'h00;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h1c;
    mem[243] = 8'h00;
    mem[244] = 8'h00;
    mem[245] = 8'h00;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'h00;
    mem[251] = 8'h00;
    mem[252] = 8'h00;
    mem[253] = 8'h00;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'h00;
    mem[259] = 8'h00;
    mem[260] = 8'h00;
    mem[261] = 8'h00;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'h00;
    mem[267] = 8'h00;
    mem[268] = 8'h00;
    mem[269] = 8'h00;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'h00;
    mem[275] = 8'h00;
    mem[276] = 8'h00;
    mem[277] = 8'h00;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h00;
    mem[283] = 8'h00;
    mem[284] = 8'h00;
    mem[285] = 8'h00;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'h00;
    mem[291] = 8'h00;
    mem[292] = 8'h00;
    mem[293] = 8'h00;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'h00;
    mem[300] = 8'h00;
    mem[301] = 8'h00;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'h00;
    mem[307] = 8'h00;
    mem[308] = 8'h00;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'h00;
    mem[316] = 8'h00;
    mem[317] = 8'h00;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'h00;
    mem[323] = 8'h00;
    mem[324] = 8'h00;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'h00;
    mem[332] = 8'h00;
    mem[333] = 8'h00;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'h00;
    mem[339] = 8'h00;
    mem[340] = 8'h00;
    mem[341] = 8'h00;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'h00;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'hfe;
    mem[354] = 8'hff;
    mem[355] = 8'hff;
    mem[356] = 8'hff;
    mem[357] = 8'hff;
    mem[358] = 8'hff;
    mem[359] = 8'h0f;
    mem[360] = 8'hf8;
    mem[361] = 8'hff;
    mem[362] = 8'hff;
    mem[363] = 8'hff;
    mem[364] = 8'hff;
    mem[365] = 8'hff;
    mem[366] = 8'h1f;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'hfe;
    mem[370] = 8'hff;
    mem[371] = 8'hff;
    mem[372] = 8'hff;
    mem[373] = 8'hff;
    mem[374] = 8'hff;
    mem[375] = 8'h1f;
    mem[376] = 8'hf8;
    mem[377] = 8'hff;
    mem[378] = 8'hff;
    mem[379] = 8'hff;
    mem[380] = 8'hff;
    mem[381] = 8'hff;
    mem[382] = 8'h1f;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'hfe;
    mem[386] = 8'hff;
    mem[387] = 8'hff;
    mem[388] = 8'hff;
    mem[389] = 8'hff;
    mem[390] = 8'hff;
    mem[391] = 8'h1f;
    mem[392] = 8'hf8;
    mem[393] = 8'hff;
    mem[394] = 8'hff;
    mem[395] = 8'hff;
    mem[396] = 8'hff;
    mem[397] = 8'hff;
    mem[398] = 8'h1f;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'hfe;
    mem[402] = 8'hff;
    mem[403] = 8'hff;
    mem[404] = 8'hff;
    mem[405] = 8'hff;
    mem[406] = 8'hff;
    mem[407] = 8'h1f;
    mem[408] = 8'hfc;
    mem[409] = 8'hff;
    mem[410] = 8'hff;
    mem[411] = 8'hff;
    mem[412] = 8'hff;
    mem[413] = 8'hff;
    mem[414] = 8'h1f;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'hfe;
    mem[418] = 8'hff;
    mem[419] = 8'hff;
    mem[420] = 8'hff;
    mem[421] = 8'hff;
    mem[422] = 8'hff;
    mem[423] = 8'h1f;
    mem[424] = 8'hf8;
    mem[425] = 8'hff;
    mem[426] = 8'hff;
    mem[427] = 8'hff;
    mem[428] = 8'hff;
    mem[429] = 8'hff;
    mem[430] = 8'h1f;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'hfe;
    mem[434] = 8'hff;
    mem[435] = 8'hff;
    mem[436] = 8'hff;
    mem[437] = 8'hff;
    mem[438] = 8'hff;
    mem[439] = 8'h1f;
    mem[440] = 8'hfc;
    mem[441] = 8'hff;
    mem[442] = 8'hff;
    mem[443] = 8'hff;
    mem[444] = 8'hff;
    mem[445] = 8'hff;
    mem[446] = 8'h1f;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'hfe;
    mem[450] = 8'hff;
    mem[451] = 8'hff;
    mem[452] = 8'hff;
    mem[453] = 8'hff;
    mem[454] = 8'hff;
    mem[455] = 8'h1f;
    mem[456] = 8'hf8;
    mem[457] = 8'hff;
    mem[458] = 8'hff;
    mem[459] = 8'hff;
    mem[460] = 8'hff;
    mem[461] = 8'hff;
    mem[462] = 8'h1f;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'hfe;
    mem[466] = 8'hff;
    mem[467] = 8'hff;
    mem[468] = 8'hff;
    mem[469] = 8'hff;
    mem[470] = 8'hff;
    mem[471] = 8'h1f;
    mem[472] = 8'hf8;
    mem[473] = 8'hff;
    mem[474] = 8'hff;
    mem[475] = 8'hff;
    mem[476] = 8'hff;
    mem[477] = 8'hff;
    mem[478] = 8'h1f;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'hfe;
    mem[482] = 8'hff;
    mem[483] = 8'hff;
    mem[484] = 8'hff;
    mem[485] = 8'hff;
    mem[486] = 8'hff;
    mem[487] = 8'h1f;
    mem[488] = 8'hf8;
    mem[489] = 8'hff;
    mem[490] = 8'hff;
    mem[491] = 8'hff;
    mem[492] = 8'hff;
    mem[493] = 8'hff;
    mem[494] = 8'h1f;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'hfe;
    mem[498] = 8'hff;
    mem[499] = 8'hff;
    mem[500] = 8'hff;
    mem[501] = 8'hff;
    mem[502] = 8'hff;
    mem[503] = 8'h1f;
    mem[504] = 8'hf8;
    mem[505] = 8'hff;
    mem[506] = 8'hff;
    mem[507] = 8'hff;
    mem[508] = 8'hff;
    mem[509] = 8'hff;
    mem[510] = 8'h1f;
    mem[511] = 8'h00;
    mem[512] = 8'h00;
    mem[513] = 8'hfe;
    mem[514] = 8'hff;
    mem[515] = 8'hff;
    mem[516] = 8'hff;
    mem[517] = 8'hff;
    mem[518] = 8'hff;
    mem[519] = 8'h1f;
    mem[520] = 8'hfc;
    mem[521] = 8'hff;
    mem[522] = 8'hff;
    mem[523] = 8'hff;
    mem[524] = 8'hff;
    mem[525] = 8'hff;
    mem[526] = 8'h1f;
    mem[527] = 8'h00;
    mem[528] = 8'h00;
    mem[529] = 8'hfe;
    mem[530] = 8'hff;
    mem[531] = 8'hff;
    mem[532] = 8'hff;
    mem[533] = 8'hff;
    mem[534] = 8'hff;
    mem[535] = 8'h1f;
    mem[536] = 8'hf8;
    mem[537] = 8'hff;
    mem[538] = 8'hff;
    mem[539] = 8'hff;
    mem[540] = 8'hff;
    mem[541] = 8'hff;
    mem[542] = 8'h1f;
    mem[543] = 8'h00;
    mem[544] = 8'h00;
    mem[545] = 8'hfe;
    mem[546] = 8'hff;
    mem[547] = 8'h07;
    mem[548] = 8'hf8;
    mem[549] = 8'hff;
    mem[550] = 8'hff;
    mem[551] = 8'h1f;
    mem[552] = 8'hfc;
    mem[553] = 8'hff;
    mem[554] = 8'hff;
    mem[555] = 8'h03;
    mem[556] = 8'he0;
    mem[557] = 8'hff;
    mem[558] = 8'h1f;
    mem[559] = 8'h00;
    mem[560] = 8'h00;
    mem[561] = 8'hfe;
    mem[562] = 8'h7f;
    mem[563] = 8'h00;
    mem[564] = 8'hc0;
    mem[565] = 8'hff;
    mem[566] = 8'hff;
    mem[567] = 8'h1f;
    mem[568] = 8'hf8;
    mem[569] = 8'hff;
    mem[570] = 8'hff;
    mem[571] = 8'h00;
    mem[572] = 8'h00;
    mem[573] = 8'hff;
    mem[574] = 8'h1f;
    mem[575] = 8'h00;
    mem[576] = 8'h00;
    mem[577] = 8'hfe;
    mem[578] = 8'h1f;
    mem[579] = 8'h00;
    mem[580] = 8'h80;
    mem[581] = 8'hff;
    mem[582] = 8'hff;
    mem[583] = 8'h1f;
    mem[584] = 8'hfc;
    mem[585] = 8'hff;
    mem[586] = 8'h7f;
    mem[587] = 8'h00;
    mem[588] = 8'h00;
    mem[589] = 8'hfe;
    mem[590] = 8'h1f;
    mem[591] = 8'h00;
    mem[592] = 8'h00;
    mem[593] = 8'hfe;
    mem[594] = 8'h1f;
    mem[595] = 8'hfc;
    mem[596] = 8'h00;
    mem[597] = 8'hff;
    mem[598] = 8'hff;
    mem[599] = 8'h1f;
    mem[600] = 8'hf8;
    mem[601] = 8'hff;
    mem[602] = 8'h3f;
    mem[603] = 8'h00;
    mem[604] = 8'h0f;
    mem[605] = 8'hfc;
    mem[606] = 8'h1f;
    mem[607] = 8'h00;
    mem[608] = 8'h00;
    mem[609] = 8'hfe;
    mem[610] = 8'h1f;
    mem[611] = 8'hff;
    mem[612] = 8'h03;
    mem[613] = 8'hfe;
    mem[614] = 8'hff;
    mem[615] = 8'h1f;
    mem[616] = 8'hf8;
    mem[617] = 8'hff;
    mem[618] = 8'h1f;
    mem[619] = 8'he0;
    mem[620] = 8'h3f;
    mem[621] = 8'hfc;
    mem[622] = 8'h1f;
    mem[623] = 8'h00;
    mem[624] = 8'h00;
    mem[625] = 8'hfe;
    mem[626] = 8'hdf;
    mem[627] = 8'hff;
    mem[628] = 8'h0f;
    mem[629] = 8'hfe;
    mem[630] = 8'hff;
    mem[631] = 8'h1f;
    mem[632] = 8'hf8;
    mem[633] = 8'hff;
    mem[634] = 8'h1f;
    mem[635] = 8'hf8;
    mem[636] = 8'hff;
    mem[637] = 8'hf8;
    mem[638] = 8'h1f;
    mem[639] = 8'h00;
    mem[640] = 8'h00;
    mem[641] = 8'hfe;
    mem[642] = 8'hff;
    mem[643] = 8'hff;
    mem[644] = 8'h0f;
    mem[645] = 8'hfe;
    mem[646] = 8'hff;
    mem[647] = 8'h1f;
    mem[648] = 8'hf8;
    mem[649] = 8'hff;
    mem[650] = 8'h1f;
    mem[651] = 8'hf8;
    mem[652] = 8'hff;
    mem[653] = 8'hf8;
    mem[654] = 8'h3f;
    mem[655] = 8'h00;
    mem[656] = 8'h00;
    mem[657] = 8'hfe;
    mem[658] = 8'hff;
    mem[659] = 8'hff;
    mem[660] = 8'h0f;
    mem[661] = 8'hfe;
    mem[662] = 8'hff;
    mem[663] = 8'h1f;
    mem[664] = 8'hfc;
    mem[665] = 8'hff;
    mem[666] = 8'h0f;
    mem[667] = 8'hfc;
    mem[668] = 8'hff;
    mem[669] = 8'hfd;
    mem[670] = 8'h1f;
    mem[671] = 8'h00;
    mem[672] = 8'h00;
    mem[673] = 8'hfe;
    mem[674] = 8'hff;
    mem[675] = 8'hff;
    mem[676] = 8'h0f;
    mem[677] = 8'hfe;
    mem[678] = 8'hff;
    mem[679] = 8'h1f;
    mem[680] = 8'hf8;
    mem[681] = 8'hff;
    mem[682] = 8'h0f;
    mem[683] = 8'hf8;
    mem[684] = 8'hff;
    mem[685] = 8'hff;
    mem[686] = 8'h1f;
    mem[687] = 8'h00;
    mem[688] = 8'h00;
    mem[689] = 8'hfe;
    mem[690] = 8'hff;
    mem[691] = 8'hff;
    mem[692] = 8'h0f;
    mem[693] = 8'hfe;
    mem[694] = 8'hff;
    mem[695] = 8'h1f;
    mem[696] = 8'hfc;
    mem[697] = 8'hff;
    mem[698] = 8'h1f;
    mem[699] = 8'hf8;
    mem[700] = 8'hff;
    mem[701] = 8'hff;
    mem[702] = 8'h3f;
    mem[703] = 8'h00;
    mem[704] = 8'h00;
    mem[705] = 8'hfe;
    mem[706] = 8'hff;
    mem[707] = 8'hff;
    mem[708] = 8'h0f;
    mem[709] = 8'hfe;
    mem[710] = 8'hff;
    mem[711] = 8'h1f;
    mem[712] = 8'hf8;
    mem[713] = 8'hff;
    mem[714] = 8'h1f;
    mem[715] = 8'hf8;
    mem[716] = 8'hff;
    mem[717] = 8'hff;
    mem[718] = 8'h3f;
    mem[719] = 8'h00;
    mem[720] = 8'h00;
    mem[721] = 8'hfe;
    mem[722] = 8'hff;
    mem[723] = 8'hff;
    mem[724] = 8'h0f;
    mem[725] = 8'hfe;
    mem[726] = 8'hff;
    mem[727] = 8'h1f;
    mem[728] = 8'hfc;
    mem[729] = 8'hff;
    mem[730] = 8'h1f;
    mem[731] = 8'hf0;
    mem[732] = 8'hff;
    mem[733] = 8'hff;
    mem[734] = 8'h3f;
    mem[735] = 8'h00;
    mem[736] = 8'h00;
    mem[737] = 8'hfe;
    mem[738] = 8'hff;
    mem[739] = 8'hff;
    mem[740] = 8'h07;
    mem[741] = 8'hfe;
    mem[742] = 8'hff;
    mem[743] = 8'h1f;
    mem[744] = 8'hfc;
    mem[745] = 8'hff;
    mem[746] = 8'h1f;
    mem[747] = 8'hf0;
    mem[748] = 8'hff;
    mem[749] = 8'hff;
    mem[750] = 8'h3f;
    mem[751] = 8'h00;
    mem[752] = 8'h00;
    mem[753] = 8'hfe;
    mem[754] = 8'hff;
    mem[755] = 8'hff;
    mem[756] = 8'h03;
    mem[757] = 8'hff;
    mem[758] = 8'hff;
    mem[759] = 8'h1f;
    mem[760] = 8'hfc;
    mem[761] = 8'hff;
    mem[762] = 8'h3f;
    mem[763] = 8'he0;
    mem[764] = 8'hff;
    mem[765] = 8'hff;
    mem[766] = 8'h3f;
    mem[767] = 8'h00;
    mem[768] = 8'h00;
    mem[769] = 8'hfe;
    mem[770] = 8'hff;
    mem[771] = 8'hff;
    mem[772] = 8'h01;
    mem[773] = 8'hff;
    mem[774] = 8'hff;
    mem[775] = 8'h1f;
    mem[776] = 8'hfc;
    mem[777] = 8'hff;
    mem[778] = 8'h3f;
    mem[779] = 8'hc0;
    mem[780] = 8'hff;
    mem[781] = 8'hff;
    mem[782] = 8'h3f;
    mem[783] = 8'h00;
    mem[784] = 8'h00;
    mem[785] = 8'hfe;
    mem[786] = 8'hff;
    mem[787] = 8'hff;
    mem[788] = 8'h80;
    mem[789] = 8'hff;
    mem[790] = 8'hff;
    mem[791] = 8'h1f;
    mem[792] = 8'hfc;
    mem[793] = 8'hff;
    mem[794] = 8'h7f;
    mem[795] = 8'h80;
    mem[796] = 8'hff;
    mem[797] = 8'hff;
    mem[798] = 8'h3f;
    mem[799] = 8'h00;
    mem[800] = 8'h00;
    mem[801] = 8'hfe;
    mem[802] = 8'hff;
    mem[803] = 8'h7f;
    mem[804] = 8'h80;
    mem[805] = 8'hff;
    mem[806] = 8'hff;
    mem[807] = 8'h1f;
    mem[808] = 8'hfc;
    mem[809] = 8'hff;
    mem[810] = 8'h7f;
    mem[811] = 8'h00;
    mem[812] = 8'hff;
    mem[813] = 8'hff;
    mem[814] = 8'h3f;
    mem[815] = 8'h00;
    mem[816] = 8'h00;
    mem[817] = 8'hfe;
    mem[818] = 8'hff;
    mem[819] = 8'h3f;
    mem[820] = 8'hc0;
    mem[821] = 8'hff;
    mem[822] = 8'hff;
    mem[823] = 8'h1f;
    mem[824] = 8'hf8;
    mem[825] = 8'hff;
    mem[826] = 8'hff;
    mem[827] = 8'h01;
    mem[828] = 8'hfe;
    mem[829] = 8'hff;
    mem[830] = 8'h3f;
    mem[831] = 8'h00;
    mem[832] = 8'h00;
    mem[833] = 8'hfe;
    mem[834] = 8'hff;
    mem[835] = 8'h1f;
    mem[836] = 8'he0;
    mem[837] = 8'hff;
    mem[838] = 8'hff;
    mem[839] = 8'h1f;
    mem[840] = 8'hfc;
    mem[841] = 8'hff;
    mem[842] = 8'hff;
    mem[843] = 8'h01;
    mem[844] = 8'hfc;
    mem[845] = 8'hff;
    mem[846] = 8'h3f;
    mem[847] = 8'h00;
    mem[848] = 8'h00;
    mem[849] = 8'hfe;
    mem[850] = 8'hff;
    mem[851] = 8'h07;
    mem[852] = 8'hf0;
    mem[853] = 8'hff;
    mem[854] = 8'hff;
    mem[855] = 8'h1f;
    mem[856] = 8'hf8;
    mem[857] = 8'hff;
    mem[858] = 8'hff;
    mem[859] = 8'h03;
    mem[860] = 8'hf0;
    mem[861] = 8'hff;
    mem[862] = 8'h3f;
    mem[863] = 8'h00;
    mem[864] = 8'h00;
    mem[865] = 8'hff;
    mem[866] = 8'hff;
    mem[867] = 8'h03;
    mem[868] = 8'hf0;
    mem[869] = 8'hff;
    mem[870] = 8'hff;
    mem[871] = 8'h1f;
    mem[872] = 8'hfc;
    mem[873] = 8'hff;
    mem[874] = 8'hff;
    mem[875] = 8'h03;
    mem[876] = 8'he0;
    mem[877] = 8'hff;
    mem[878] = 8'h3f;
    mem[879] = 8'h00;
    mem[880] = 8'h00;
    mem[881] = 8'hff;
    mem[882] = 8'hff;
    mem[883] = 8'h01;
    mem[884] = 8'hf8;
    mem[885] = 8'hff;
    mem[886] = 8'hff;
    mem[887] = 8'h1f;
    mem[888] = 8'hf8;
    mem[889] = 8'hff;
    mem[890] = 8'hff;
    mem[891] = 8'h0f;
    mem[892] = 8'hc0;
    mem[893] = 8'hff;
    mem[894] = 8'h3f;
    mem[895] = 8'h00;
    mem[896] = 8'h00;
    mem[897] = 8'hff;
    mem[898] = 8'hff;
    mem[899] = 8'h00;
    mem[900] = 8'hfc;
    mem[901] = 8'hff;
    mem[902] = 8'hff;
    mem[903] = 8'h1f;
    mem[904] = 8'hf8;
    mem[905] = 8'hff;
    mem[906] = 8'hff;
    mem[907] = 8'h0f;
    mem[908] = 8'h00;
    mem[909] = 8'hff;
    mem[910] = 8'h3f;
    mem[911] = 8'h00;
    mem[912] = 8'h00;
    mem[913] = 8'hff;
    mem[914] = 8'h1f;
    mem[915] = 8'h00;
    mem[916] = 8'hff;
    mem[917] = 8'hff;
    mem[918] = 8'hff;
    mem[919] = 8'h1f;
    mem[920] = 8'hf8;
    mem[921] = 8'hff;
    mem[922] = 8'hff;
    mem[923] = 8'h1f;
    mem[924] = 8'h00;
    mem[925] = 8'hfe;
    mem[926] = 8'h3f;
    mem[927] = 8'h00;
    mem[928] = 8'h00;
    mem[929] = 8'hff;
    mem[930] = 8'h1f;
    mem[931] = 8'h00;
    mem[932] = 8'hff;
    mem[933] = 8'hff;
    mem[934] = 8'hff;
    mem[935] = 8'h1f;
    mem[936] = 8'hfc;
    mem[937] = 8'hff;
    mem[938] = 8'hff;
    mem[939] = 8'h3f;
    mem[940] = 8'h00;
    mem[941] = 8'hf8;
    mem[942] = 8'h3f;
    mem[943] = 8'h00;
    mem[944] = 8'h00;
    mem[945] = 8'hff;
    mem[946] = 8'h07;
    mem[947] = 8'h80;
    mem[948] = 8'hff;
    mem[949] = 8'hff;
    mem[950] = 8'hff;
    mem[951] = 8'h1f;
    mem[952] = 8'hfc;
    mem[953] = 8'hff;
    mem[954] = 8'hff;
    mem[955] = 8'h7f;
    mem[956] = 8'h00;
    mem[957] = 8'hf8;
    mem[958] = 8'h3f;
    mem[959] = 8'h00;
    mem[960] = 8'h00;
    mem[961] = 8'hff;
    mem[962] = 8'h03;
    mem[963] = 8'hc0;
    mem[964] = 8'hff;
    mem[965] = 8'hff;
    mem[966] = 8'hff;
    mem[967] = 8'h1f;
    mem[968] = 8'hf8;
    mem[969] = 8'hff;
    mem[970] = 8'hff;
    mem[971] = 8'hff;
    mem[972] = 8'h00;
    mem[973] = 8'hc0;
    mem[974] = 8'h3f;
    mem[975] = 8'h00;
    mem[976] = 8'h00;
    mem[977] = 8'hff;
    mem[978] = 8'h00;
    mem[979] = 8'hf0;
    mem[980] = 8'hff;
    mem[981] = 8'hff;
    mem[982] = 8'hff;
    mem[983] = 8'h0f;
    mem[984] = 8'hf8;
    mem[985] = 8'hff;
    mem[986] = 8'hff;
    mem[987] = 8'hff;
    mem[988] = 8'h01;
    mem[989] = 8'h80;
    mem[990] = 8'h3f;
    mem[991] = 8'h00;
    mem[992] = 8'h00;
    mem[993] = 8'h3f;
    mem[994] = 8'h00;
    mem[995] = 8'hf0;
    mem[996] = 8'hff;
    mem[997] = 8'hff;
    mem[998] = 8'hff;
    mem[999] = 8'h0f;
    mem[1000] = 8'hf0;
    mem[1001] = 8'hff;
    mem[1002] = 8'hff;
    mem[1003] = 8'hff;
    mem[1004] = 8'h03;
    mem[1005] = 8'h00;
    mem[1006] = 8'h3e;
    mem[1007] = 8'h00;
    mem[1008] = 8'h00;
    mem[1009] = 8'h1f;
    mem[1010] = 8'h00;
    mem[1011] = 8'hf8;
    mem[1012] = 8'hff;
    mem[1013] = 8'hff;
    mem[1014] = 8'hff;
    mem[1015] = 8'h03;
    mem[1016] = 8'hc0;
    mem[1017] = 8'hff;
    mem[1018] = 8'hff;
    mem[1019] = 8'hff;
    mem[1020] = 8'h0f;
    mem[1021] = 8'h00;
    mem[1022] = 8'h38;
    mem[1023] = 8'h00;
    mem[1024] = 8'h00;
    mem[1025] = 8'h07;
    mem[1026] = 8'h00;
    mem[1027] = 8'hfe;
    mem[1028] = 8'hff;
    mem[1029] = 8'hff;
    mem[1030] = 8'hff;
    mem[1031] = 8'h00;
    mem[1032] = 8'h80;
    mem[1033] = 8'hff;
    mem[1034] = 8'hff;
    mem[1035] = 8'hff;
    mem[1036] = 8'h1f;
    mem[1037] = 8'h00;
    mem[1038] = 8'h30;
    mem[1039] = 8'h00;
    mem[1040] = 8'h00;
    mem[1041] = 8'h03;
    mem[1042] = 8'h00;
    mem[1043] = 8'hfe;
    mem[1044] = 8'hff;
    mem[1045] = 8'hff;
    mem[1046] = 8'h7f;
    mem[1047] = 8'h00;
    mem[1048] = 8'h00;
    mem[1049] = 8'hff;
    mem[1050] = 8'hff;
    mem[1051] = 8'hff;
    mem[1052] = 8'h1f;
    mem[1053] = 8'h00;
    mem[1054] = 8'h30;
    mem[1055] = 8'h00;
    mem[1056] = 8'h00;
    mem[1057] = 8'h03;
    mem[1058] = 8'h00;
    mem[1059] = 8'hff;
    mem[1060] = 8'hff;
    mem[1061] = 8'hff;
    mem[1062] = 8'h1f;
    mem[1063] = 8'h00;
    mem[1064] = 8'h00;
    mem[1065] = 8'hfe;
    mem[1066] = 8'hff;
    mem[1067] = 8'hff;
    mem[1068] = 8'h3f;
    mem[1069] = 8'h00;
    mem[1070] = 8'h20;
    mem[1071] = 8'h00;
    mem[1072] = 8'h00;
    mem[1073] = 8'h03;
    mem[1074] = 8'h80;
    mem[1075] = 8'hff;
    mem[1076] = 8'hff;
    mem[1077] = 8'hff;
    mem[1078] = 8'h0f;
    mem[1079] = 8'h00;
    mem[1080] = 8'h00;
    mem[1081] = 8'hf8;
    mem[1082] = 8'hff;
    mem[1083] = 8'hff;
    mem[1084] = 8'h7f;
    mem[1085] = 8'h00;
    mem[1086] = 8'h00;
    mem[1087] = 8'h00;
    mem[1088] = 8'h00;
    mem[1089] = 8'h00;
    mem[1090] = 8'hc0;
    mem[1091] = 8'hff;
    mem[1092] = 8'hff;
    mem[1093] = 8'hff;
    mem[1094] = 8'h07;
    mem[1095] = 8'h00;
    mem[1096] = 8'h00;
    mem[1097] = 8'hf0;
    mem[1098] = 8'hff;
    mem[1099] = 8'hff;
    mem[1100] = 8'hff;
    mem[1101] = 8'h00;
    mem[1102] = 8'h00;
    mem[1103] = 8'h00;
    mem[1104] = 8'h00;
    mem[1105] = 8'h00;
    mem[1106] = 8'he0;
    mem[1107] = 8'hff;
    mem[1108] = 8'hff;
    mem[1109] = 8'hff;
    mem[1110] = 8'h03;
    mem[1111] = 8'h00;
    mem[1112] = 8'h00;
    mem[1113] = 8'he0;
    mem[1114] = 8'hff;
    mem[1115] = 8'hff;
    mem[1116] = 8'hff;
    mem[1117] = 8'h01;
    mem[1118] = 8'h00;
    mem[1119] = 8'h00;
    mem[1120] = 8'h00;
    mem[1121] = 8'h00;
    mem[1122] = 8'he0;
    mem[1123] = 8'hff;
    mem[1124] = 8'hff;
    mem[1125] = 8'hff;
    mem[1126] = 8'h01;
    mem[1127] = 8'h00;
    mem[1128] = 8'h00;
    mem[1129] = 8'hc0;
    mem[1130] = 8'hff;
    mem[1131] = 8'hff;
    mem[1132] = 8'hff;
    mem[1133] = 8'h01;
    mem[1134] = 8'h00;
    mem[1135] = 8'h00;
    mem[1136] = 8'h00;
    mem[1137] = 8'h00;
    mem[1138] = 8'hf0;
    mem[1139] = 8'hff;
    mem[1140] = 8'hff;
    mem[1141] = 8'hff;
    mem[1142] = 8'h00;
    mem[1143] = 8'h00;
    mem[1144] = 8'h00;
    mem[1145] = 8'h80;
    mem[1146] = 8'hff;
    mem[1147] = 8'hff;
    mem[1148] = 8'hff;
    mem[1149] = 8'h03;
    mem[1150] = 8'h00;
    mem[1151] = 8'h00;
    mem[1152] = 8'h00;
    mem[1153] = 8'h00;
    mem[1154] = 8'hf8;
    mem[1155] = 8'hff;
    mem[1156] = 8'hff;
    mem[1157] = 8'h7f;
    mem[1158] = 8'h00;
    mem[1159] = 8'h00;
    mem[1160] = 8'h00;
    mem[1161] = 8'h00;
    mem[1162] = 8'hff;
    mem[1163] = 8'hff;
    mem[1164] = 8'hff;
    mem[1165] = 8'h07;
    mem[1166] = 8'h00;
    mem[1167] = 8'h00;
    mem[1168] = 8'h00;
    mem[1169] = 8'h00;
    mem[1170] = 8'hf8;
    mem[1171] = 8'hff;
    mem[1172] = 8'hff;
    mem[1173] = 8'h3f;
    mem[1174] = 8'h00;
    mem[1175] = 8'h00;
    mem[1176] = 8'h00;
    mem[1177] = 8'h00;
    mem[1178] = 8'hfe;
    mem[1179] = 8'hff;
    mem[1180] = 8'hff;
    mem[1181] = 8'h07;
    mem[1182] = 8'h00;
    mem[1183] = 8'h00;
    mem[1184] = 8'h00;
    mem[1185] = 8'h00;
    mem[1186] = 8'hfc;
    mem[1187] = 8'hff;
    mem[1188] = 8'hff;
    mem[1189] = 8'h1f;
    mem[1190] = 8'h00;
    mem[1191] = 8'h00;
    mem[1192] = 8'h00;
    mem[1193] = 8'h00;
    mem[1194] = 8'hfc;
    mem[1195] = 8'hff;
    mem[1196] = 8'hff;
    mem[1197] = 8'h07;
    mem[1198] = 8'h00;
    mem[1199] = 8'h00;
    mem[1200] = 8'h00;
    mem[1201] = 8'h00;
    mem[1202] = 8'hfc;
    mem[1203] = 8'hff;
    mem[1204] = 8'hff;
    mem[1205] = 8'h1f;
    mem[1206] = 8'h00;
    mem[1207] = 8'h00;
    mem[1208] = 8'h00;
    mem[1209] = 8'h00;
    mem[1210] = 8'hfc;
    mem[1211] = 8'hff;
    mem[1212] = 8'hff;
    mem[1213] = 8'h0f;
    mem[1214] = 8'h00;
    mem[1215] = 8'h00;
    mem[1216] = 8'h00;
    mem[1217] = 8'h00;
    mem[1218] = 8'hfc;
    mem[1219] = 8'hff;
    mem[1220] = 8'hff;
    mem[1221] = 8'h0f;
    mem[1222] = 8'h00;
    mem[1223] = 8'h00;
    mem[1224] = 8'h00;
    mem[1225] = 8'h00;
    mem[1226] = 8'hfc;
    mem[1227] = 8'hff;
    mem[1228] = 8'hff;
    mem[1229] = 8'h1f;
    mem[1230] = 8'h00;
    mem[1231] = 8'h00;
    mem[1232] = 8'h00;
    mem[1233] = 8'h00;
    mem[1234] = 8'hfc;
    mem[1235] = 8'hff;
    mem[1236] = 8'hff;
    mem[1237] = 8'h0f;
    mem[1238] = 8'h00;
    mem[1239] = 8'h00;
    mem[1240] = 8'h00;
    mem[1241] = 8'h00;
    mem[1242] = 8'hf8;
    mem[1243] = 8'hff;
    mem[1244] = 8'hff;
    mem[1245] = 8'h1f;
    mem[1246] = 8'h00;
    mem[1247] = 8'h00;
    mem[1248] = 8'h00;
    mem[1249] = 8'h00;
    mem[1250] = 8'hfe;
    mem[1251] = 8'hff;
    mem[1252] = 8'hff;
    mem[1253] = 8'h07;
    mem[1254] = 8'h00;
    mem[1255] = 8'h00;
    mem[1256] = 8'h00;
    mem[1257] = 8'h00;
    mem[1258] = 8'hf0;
    mem[1259] = 8'hff;
    mem[1260] = 8'hff;
    mem[1261] = 8'h1f;
    mem[1262] = 8'h00;
    mem[1263] = 8'h00;
    mem[1264] = 8'h00;
    mem[1265] = 8'h00;
    mem[1266] = 8'hfe;
    mem[1267] = 8'hff;
    mem[1268] = 8'hff;
    mem[1269] = 8'h07;
    mem[1270] = 8'h00;
    mem[1271] = 8'h00;
    mem[1272] = 8'h00;
    mem[1273] = 8'h00;
    mem[1274] = 8'hf0;
    mem[1275] = 8'hff;
    mem[1276] = 8'hff;
    mem[1277] = 8'h1f;
    mem[1278] = 8'h00;
    mem[1279] = 8'h00;
    mem[1280] = 8'h00;
    mem[1281] = 8'h00;
    mem[1282] = 8'hfe;
    mem[1283] = 8'hff;
    mem[1284] = 8'hff;
    mem[1285] = 8'h07;
    mem[1286] = 8'h00;
    mem[1287] = 8'h00;
    mem[1288] = 8'h00;
    mem[1289] = 8'h00;
    mem[1290] = 8'hf0;
    mem[1291] = 8'hff;
    mem[1292] = 8'hff;
    mem[1293] = 8'h1f;
    mem[1294] = 8'h00;
    mem[1295] = 8'h00;
    mem[1296] = 8'h00;
    mem[1297] = 8'h00;
    mem[1298] = 8'hfe;
    mem[1299] = 8'hff;
    mem[1300] = 8'hff;
    mem[1301] = 8'h07;
    mem[1302] = 8'h00;
    mem[1303] = 8'h00;
    mem[1304] = 8'h00;
    mem[1305] = 8'h00;
    mem[1306] = 8'hf0;
    mem[1307] = 8'hff;
    mem[1308] = 8'hff;
    mem[1309] = 8'h1f;
    mem[1310] = 8'h00;
    mem[1311] = 8'h00;
    mem[1312] = 8'h00;
    mem[1313] = 8'h00;
    mem[1314] = 8'hfe;
    mem[1315] = 8'hff;
    mem[1316] = 8'hff;
    mem[1317] = 8'h07;
    mem[1318] = 8'h00;
    mem[1319] = 8'h00;
    mem[1320] = 8'h00;
    mem[1321] = 8'h00;
    mem[1322] = 8'hf0;
    mem[1323] = 8'hff;
    mem[1324] = 8'hff;
    mem[1325] = 8'h1f;
    mem[1326] = 8'h00;
    mem[1327] = 8'h00;
    mem[1328] = 8'h00;
    mem[1329] = 8'h00;
    mem[1330] = 8'hfe;
    mem[1331] = 8'hff;
    mem[1332] = 8'hff;
    mem[1333] = 8'h07;
    mem[1334] = 8'h00;
    mem[1335] = 8'h00;
    mem[1336] = 8'h00;
    mem[1337] = 8'h00;
    mem[1338] = 8'hf0;
    mem[1339] = 8'hff;
    mem[1340] = 8'hff;
    mem[1341] = 8'h1f;
    mem[1342] = 8'h00;
    mem[1343] = 8'h00;
    mem[1344] = 8'h00;
    mem[1345] = 8'h00;
    mem[1346] = 8'hfe;
    mem[1347] = 8'hff;
    mem[1348] = 8'hff;
    mem[1349] = 8'h07;
    mem[1350] = 8'h00;
    mem[1351] = 8'h00;
    mem[1352] = 8'h00;
    mem[1353] = 8'h00;
    mem[1354] = 8'hf0;
    mem[1355] = 8'hff;
    mem[1356] = 8'hff;
    mem[1357] = 8'h1f;
    mem[1358] = 8'h00;
    mem[1359] = 8'h00;
    mem[1360] = 8'h00;
    mem[1361] = 8'h00;
    mem[1362] = 8'hfc;
    mem[1363] = 8'hff;
    mem[1364] = 8'hff;
    mem[1365] = 8'h0f;
    mem[1366] = 8'h00;
    mem[1367] = 8'h00;
    mem[1368] = 8'h00;
    mem[1369] = 8'h00;
    mem[1370] = 8'hf8;
    mem[1371] = 8'hff;
    mem[1372] = 8'hff;
    mem[1373] = 8'h1f;
    mem[1374] = 8'h00;
    mem[1375] = 8'h00;
    mem[1376] = 8'h00;
    mem[1377] = 8'h00;
    mem[1378] = 8'hfc;
    mem[1379] = 8'hff;
    mem[1380] = 8'hff;
    mem[1381] = 8'h0f;
    mem[1382] = 8'h00;
    mem[1383] = 8'h00;
    mem[1384] = 8'h00;
    mem[1385] = 8'h00;
    mem[1386] = 8'hfc;
    mem[1387] = 8'hff;
    mem[1388] = 8'hff;
    mem[1389] = 8'h1f;
    mem[1390] = 8'h00;
    mem[1391] = 8'h00;
    mem[1392] = 8'h00;
    mem[1393] = 8'h00;
    mem[1394] = 8'hfc;
    mem[1395] = 8'hff;
    mem[1396] = 8'hff;
    mem[1397] = 8'h1f;
    mem[1398] = 8'h00;
    mem[1399] = 8'h00;
    mem[1400] = 8'h00;
    mem[1401] = 8'h00;
    mem[1402] = 8'hfc;
    mem[1403] = 8'hff;
    mem[1404] = 8'hff;
    mem[1405] = 8'h0f;
    mem[1406] = 8'h00;
    mem[1407] = 8'h00;
    mem[1408] = 8'h00;
    mem[1409] = 8'h00;
    mem[1410] = 8'hfc;
    mem[1411] = 8'hff;
    mem[1412] = 8'hff;
    mem[1413] = 8'h3f;
    mem[1414] = 8'h00;
    mem[1415] = 8'h00;
    mem[1416] = 8'h00;
    mem[1417] = 8'h00;
    mem[1418] = 8'hfe;
    mem[1419] = 8'hff;
    mem[1420] = 8'hff;
    mem[1421] = 8'h07;
    mem[1422] = 8'h00;
    mem[1423] = 8'h00;
    mem[1424] = 8'h00;
    mem[1425] = 8'h00;
    mem[1426] = 8'hf8;
    mem[1427] = 8'hff;
    mem[1428] = 8'hff;
    mem[1429] = 8'h7f;
    mem[1430] = 8'h00;
    mem[1431] = 8'h00;
    mem[1432] = 8'h00;
    mem[1433] = 8'h00;
    mem[1434] = 8'hff;
    mem[1435] = 8'hff;
    mem[1436] = 8'hff;
    mem[1437] = 8'h07;
    mem[1438] = 8'h00;
    mem[1439] = 8'h00;
    mem[1440] = 8'h00;
    mem[1441] = 8'h00;
    mem[1442] = 8'hf8;
    mem[1443] = 8'hff;
    mem[1444] = 8'hff;
    mem[1445] = 8'hff;
    mem[1446] = 8'h00;
    mem[1447] = 8'h00;
    mem[1448] = 8'h00;
    mem[1449] = 8'h80;
    mem[1450] = 8'hff;
    mem[1451] = 8'hff;
    mem[1452] = 8'hff;
    mem[1453] = 8'h07;
    mem[1454] = 8'h00;
    mem[1455] = 8'h00;
    mem[1456] = 8'h00;
    mem[1457] = 8'h00;
    mem[1458] = 8'hf0;
    mem[1459] = 8'hff;
    mem[1460] = 8'hff;
    mem[1461] = 8'hff;
    mem[1462] = 8'h01;
    mem[1463] = 8'h00;
    mem[1464] = 8'h00;
    mem[1465] = 8'hc0;
    mem[1466] = 8'hff;
    mem[1467] = 8'hff;
    mem[1468] = 8'hff;
    mem[1469] = 8'h03;
    mem[1470] = 8'h00;
    mem[1471] = 8'h00;
    mem[1472] = 8'h00;
    mem[1473] = 8'h00;
    mem[1474] = 8'he0;
    mem[1475] = 8'hff;
    mem[1476] = 8'hff;
    mem[1477] = 8'hff;
    mem[1478] = 8'h03;
    mem[1479] = 8'h00;
    mem[1480] = 8'h00;
    mem[1481] = 8'hf0;
    mem[1482] = 8'hff;
    mem[1483] = 8'hff;
    mem[1484] = 8'hff;
    mem[1485] = 8'h01;
    mem[1486] = 8'h00;
    mem[1487] = 8'h00;
    mem[1488] = 8'h00;
    mem[1489] = 8'h00;
    mem[1490] = 8'he0;
    mem[1491] = 8'hff;
    mem[1492] = 8'hff;
    mem[1493] = 8'hff;
    mem[1494] = 8'h1f;
    mem[1495] = 8'h00;
    mem[1496] = 8'h00;
    mem[1497] = 8'hf8;
    mem[1498] = 8'hff;
    mem[1499] = 8'hff;
    mem[1500] = 8'hff;
    mem[1501] = 8'h00;
    mem[1502] = 8'h00;
    mem[1503] = 8'h00;
    mem[1504] = 8'h00;
    mem[1505] = 8'h00;
    mem[1506] = 8'h80;
    mem[1507] = 8'hff;
    mem[1508] = 8'hff;
    mem[1509] = 8'hff;
    mem[1510] = 8'h7f;
    mem[1511] = 8'h00;
    mem[1512] = 8'h00;
    mem[1513] = 8'hfe;
    mem[1514] = 8'hff;
    mem[1515] = 8'hff;
    mem[1516] = 8'h7f;
    mem[1517] = 8'h00;
    mem[1518] = 8'h00;
    mem[1519] = 8'h00;
    mem[1520] = 8'h00;
    mem[1521] = 8'h00;
    mem[1522] = 8'h00;
    mem[1523] = 8'hff;
    mem[1524] = 8'hff;
    mem[1525] = 8'hff;
    mem[1526] = 8'hff;
    mem[1527] = 8'h00;
    mem[1528] = 8'h80;
    mem[1529] = 8'hff;
    mem[1530] = 8'hff;
    mem[1531] = 8'hff;
    mem[1532] = 8'h7f;
    mem[1533] = 8'h00;
    mem[1534] = 8'h00;
    mem[1535] = 8'h00;
    mem[1536] = 8'h00;
    mem[1537] = 8'h00;
    mem[1538] = 8'h00;
    mem[1539] = 8'hfe;
    mem[1540] = 8'hff;
    mem[1541] = 8'hff;
    mem[1542] = 8'hff;
    mem[1543] = 8'h03;
    mem[1544] = 8'hc0;
    mem[1545] = 8'hff;
    mem[1546] = 8'hff;
    mem[1547] = 8'hff;
    mem[1548] = 8'h3f;
    mem[1549] = 8'h00;
    mem[1550] = 8'h00;
    mem[1551] = 8'h00;
    mem[1552] = 8'h00;
    mem[1553] = 8'h00;
    mem[1554] = 8'h00;
    mem[1555] = 8'hfe;
    mem[1556] = 8'hff;
    mem[1557] = 8'hff;
    mem[1558] = 8'hff;
    mem[1559] = 8'h0f;
    mem[1560] = 8'hf8;
    mem[1561] = 8'hff;
    mem[1562] = 8'hff;
    mem[1563] = 8'hff;
    mem[1564] = 8'h1f;
    mem[1565] = 8'h00;
    mem[1566] = 8'h00;
    mem[1567] = 8'h00;
    mem[1568] = 8'h00;
    mem[1569] = 8'h00;
    mem[1570] = 8'h00;
    mem[1571] = 8'hf8;
    mem[1572] = 8'hff;
    mem[1573] = 8'hff;
    mem[1574] = 8'hff;
    mem[1575] = 8'h1f;
    mem[1576] = 8'hf8;
    mem[1577] = 8'hff;
    mem[1578] = 8'hff;
    mem[1579] = 8'hff;
    mem[1580] = 8'h0f;
    mem[1581] = 8'h00;
    mem[1582] = 8'h00;
    mem[1583] = 8'h00;
    mem[1584] = 8'h00;
    mem[1585] = 8'h00;
    mem[1586] = 8'h00;
    mem[1587] = 8'hf0;
    mem[1588] = 8'hff;
    mem[1589] = 8'hff;
    mem[1590] = 8'hff;
    mem[1591] = 8'h1f;
    mem[1592] = 8'hfc;
    mem[1593] = 8'hff;
    mem[1594] = 8'hff;
    mem[1595] = 8'hff;
    mem[1596] = 8'h03;
    mem[1597] = 8'h00;
    mem[1598] = 8'h00;
    mem[1599] = 8'h00;
    mem[1600] = 8'h00;
    mem[1601] = 8'h00;
    mem[1602] = 8'h00;
    mem[1603] = 8'hc0;
    mem[1604] = 8'hff;
    mem[1605] = 8'hff;
    mem[1606] = 8'hff;
    mem[1607] = 8'h1f;
    mem[1608] = 8'hfc;
    mem[1609] = 8'hff;
    mem[1610] = 8'hff;
    mem[1611] = 8'hff;
    mem[1612] = 8'h00;
    mem[1613] = 8'h00;
    mem[1614] = 8'h00;
    mem[1615] = 8'h00;
    mem[1616] = 8'h00;
    mem[1617] = 8'h00;
    mem[1618] = 8'h00;
    mem[1619] = 8'hc0;
    mem[1620] = 8'hff;
    mem[1621] = 8'hff;
    mem[1622] = 8'hff;
    mem[1623] = 8'h1f;
    mem[1624] = 8'hfc;
    mem[1625] = 8'hff;
    mem[1626] = 8'hff;
    mem[1627] = 8'hff;
    mem[1628] = 8'h00;
    mem[1629] = 8'h00;
    mem[1630] = 8'h00;
    mem[1631] = 8'h00;
    mem[1632] = 8'h00;
    mem[1633] = 8'h00;
    mem[1634] = 8'h00;
    mem[1635] = 8'h00;
    mem[1636] = 8'hff;
    mem[1637] = 8'hff;
    mem[1638] = 8'hff;
    mem[1639] = 8'h1f;
    mem[1640] = 8'hf8;
    mem[1641] = 8'hff;
    mem[1642] = 8'hff;
    mem[1643] = 8'h7f;
    mem[1644] = 8'h00;
    mem[1645] = 8'h00;
    mem[1646] = 8'h00;
    mem[1647] = 8'h00;
    mem[1648] = 8'h00;
    mem[1649] = 8'h00;
    mem[1650] = 8'h00;
    mem[1651] = 8'h00;
    mem[1652] = 8'hfe;
    mem[1653] = 8'hff;
    mem[1654] = 8'hff;
    mem[1655] = 8'h1f;
    mem[1656] = 8'hfc;
    mem[1657] = 8'hff;
    mem[1658] = 8'hff;
    mem[1659] = 8'h1f;
    mem[1660] = 8'h00;
    mem[1661] = 8'h00;
    mem[1662] = 8'h00;
    mem[1663] = 8'h00;
    mem[1664] = 8'h00;
    mem[1665] = 8'h00;
    mem[1666] = 8'h00;
    mem[1667] = 8'h00;
    mem[1668] = 8'hf8;
    mem[1669] = 8'hff;
    mem[1670] = 8'hff;
    mem[1671] = 8'h1f;
    mem[1672] = 8'hfc;
    mem[1673] = 8'hff;
    mem[1674] = 8'hff;
    mem[1675] = 8'h07;
    mem[1676] = 8'h00;
    mem[1677] = 8'h00;
    mem[1678] = 8'h00;
    mem[1679] = 8'h00;
    mem[1680] = 8'h00;
    mem[1681] = 8'h00;
    mem[1682] = 8'h00;
    mem[1683] = 8'h00;
    mem[1684] = 8'hf0;
    mem[1685] = 8'hff;
    mem[1686] = 8'hff;
    mem[1687] = 8'h1f;
    mem[1688] = 8'hf8;
    mem[1689] = 8'hff;
    mem[1690] = 8'hff;
    mem[1691] = 8'h03;
    mem[1692] = 8'h00;
    mem[1693] = 8'h00;
    mem[1694] = 8'h00;
    mem[1695] = 8'h00;
    mem[1696] = 8'h00;
    mem[1697] = 8'h00;
    mem[1698] = 8'h00;
    mem[1699] = 8'h00;
    mem[1700] = 8'hc0;
    mem[1701] = 8'hff;
    mem[1702] = 8'hff;
    mem[1703] = 8'h1f;
    mem[1704] = 8'hfc;
    mem[1705] = 8'hff;
    mem[1706] = 8'hff;
    mem[1707] = 8'h00;
    mem[1708] = 8'h00;
    mem[1709] = 8'h00;
    mem[1710] = 8'h00;
    mem[1711] = 8'h00;
    mem[1712] = 8'h00;
    mem[1713] = 8'h00;
    mem[1714] = 8'h00;
    mem[1715] = 8'h00;
    mem[1716] = 8'h80;
    mem[1717] = 8'hff;
    mem[1718] = 8'hff;
    mem[1719] = 8'h1f;
    mem[1720] = 8'hf8;
    mem[1721] = 8'hff;
    mem[1722] = 8'h7f;
    mem[1723] = 8'h00;
    mem[1724] = 8'h00;
    mem[1725] = 8'h00;
    mem[1726] = 8'h00;
    mem[1727] = 8'h00;
    mem[1728] = 8'h00;
    mem[1729] = 8'h00;
    mem[1730] = 8'h00;
    mem[1731] = 8'h00;
    mem[1732] = 8'h00;
    mem[1733] = 8'hff;
    mem[1734] = 8'hff;
    mem[1735] = 8'h1f;
    mem[1736] = 8'hfc;
    mem[1737] = 8'hff;
    mem[1738] = 8'h1f;
    mem[1739] = 8'h00;
    mem[1740] = 8'h00;
    mem[1741] = 8'h00;
    mem[1742] = 8'h00;
    mem[1743] = 8'h00;
    mem[1744] = 8'h00;
    mem[1745] = 8'h00;
    mem[1746] = 8'h00;
    mem[1747] = 8'h00;
    mem[1748] = 8'h00;
    mem[1749] = 8'hf8;
    mem[1750] = 8'hff;
    mem[1751] = 8'h1f;
    mem[1752] = 8'hf8;
    mem[1753] = 8'hff;
    mem[1754] = 8'h07;
    mem[1755] = 8'h00;
    mem[1756] = 8'h00;
    mem[1757] = 8'h00;
    mem[1758] = 8'h00;
    mem[1759] = 8'h00;
    mem[1760] = 8'h00;
    mem[1761] = 8'h00;
    mem[1762] = 8'h00;
    mem[1763] = 8'h00;
    mem[1764] = 8'h00;
    mem[1765] = 8'hf0;
    mem[1766] = 8'hff;
    mem[1767] = 8'h1f;
    mem[1768] = 8'hf8;
    mem[1769] = 8'hff;
    mem[1770] = 8'h03;
    mem[1771] = 8'h00;
    mem[1772] = 8'h00;
    mem[1773] = 8'h00;
    mem[1774] = 8'h00;
    mem[1775] = 8'h00;
    mem[1776] = 8'h00;
    mem[1777] = 8'h00;
    mem[1778] = 8'h00;
    mem[1779] = 8'h00;
    mem[1780] = 8'h00;
    mem[1781] = 8'hc0;
    mem[1782] = 8'hff;
    mem[1783] = 8'h1f;
    mem[1784] = 8'hf8;
    mem[1785] = 8'hff;
    mem[1786] = 8'h01;
    mem[1787] = 8'h00;
    mem[1788] = 8'h00;
    mem[1789] = 8'h00;
    mem[1790] = 8'h00;
    mem[1791] = 8'h00;
    mem[1792] = 8'h00;
    mem[1793] = 8'h00;
    mem[1794] = 8'h00;
    mem[1795] = 8'h00;
    mem[1796] = 8'h00;
    mem[1797] = 8'h80;
    mem[1798] = 8'hff;
    mem[1799] = 8'h1f;
    mem[1800] = 8'hfc;
    mem[1801] = 8'h7f;
    mem[1802] = 8'h00;
    mem[1803] = 8'h00;
    mem[1804] = 8'h00;
    mem[1805] = 8'h00;
    mem[1806] = 8'h00;
    mem[1807] = 8'h00;
    mem[1808] = 8'h00;
    mem[1809] = 8'h00;
    mem[1810] = 8'h00;
    mem[1811] = 8'h00;
    mem[1812] = 8'h00;
    mem[1813] = 8'h00;
    mem[1814] = 8'hff;
    mem[1815] = 8'h1f;
    mem[1816] = 8'hf8;
    mem[1817] = 8'h3f;
    mem[1818] = 8'h00;
    mem[1819] = 8'h00;
    mem[1820] = 8'h00;
    mem[1821] = 8'h00;
    mem[1822] = 8'h00;
    mem[1823] = 8'h00;
    mem[1824] = 8'h00;
    mem[1825] = 8'h00;
    mem[1826] = 8'h00;
    mem[1827] = 8'h00;
    mem[1828] = 8'h00;
    mem[1829] = 8'h00;
    mem[1830] = 8'hfc;
    mem[1831] = 8'h1f;
    mem[1832] = 8'hf8;
    mem[1833] = 8'h0f;
    mem[1834] = 8'h00;
    mem[1835] = 8'h00;
    mem[1836] = 8'h00;
    mem[1837] = 8'h00;
    mem[1838] = 8'h00;
    mem[1839] = 8'h00;
    mem[1840] = 8'h00;
    mem[1841] = 8'h00;
    mem[1842] = 8'h00;
    mem[1843] = 8'h00;
    mem[1844] = 8'h00;
    mem[1845] = 8'h00;
    mem[1846] = 8'hf8;
    mem[1847] = 8'h1f;
    mem[1848] = 8'hfc;
    mem[1849] = 8'h07;
    mem[1850] = 8'h00;
    mem[1851] = 8'h00;
    mem[1852] = 8'h00;
    mem[1853] = 8'h00;
    mem[1854] = 8'h00;
    mem[1855] = 8'h00;
    mem[1856] = 8'h00;
    mem[1857] = 8'h00;
    mem[1858] = 8'h00;
    mem[1859] = 8'h00;
    mem[1860] = 8'h00;
    mem[1861] = 8'h00;
    mem[1862] = 8'he0;
    mem[1863] = 8'h1f;
    mem[1864] = 8'hf8;
    mem[1865] = 8'h03;
    mem[1866] = 8'h00;
    mem[1867] = 8'h00;
    mem[1868] = 8'h00;
    mem[1869] = 8'h00;
    mem[1870] = 8'h00;
    mem[1871] = 8'h00;
    mem[1872] = 8'h00;
    mem[1873] = 8'h00;
    mem[1874] = 8'h00;
    mem[1875] = 8'h00;
    mem[1876] = 8'h00;
    mem[1877] = 8'h00;
    mem[1878] = 8'he0;
    mem[1879] = 8'h1f;
    mem[1880] = 8'hfc;
    mem[1881] = 8'h00;
    mem[1882] = 8'h00;
    mem[1883] = 8'h00;
    mem[1884] = 8'h00;
    mem[1885] = 8'h00;
    mem[1886] = 8'h00;
    mem[1887] = 8'h00;
    mem[1888] = 8'h00;
    mem[1889] = 8'h00;
    mem[1890] = 8'h00;
    mem[1891] = 8'h00;
    mem[1892] = 8'h00;
    mem[1893] = 8'h00;
    mem[1894] = 8'h80;
    mem[1895] = 8'h1f;
    mem[1896] = 8'h78;
    mem[1897] = 8'h00;
    mem[1898] = 8'h00;
    mem[1899] = 8'h00;
    mem[1900] = 8'h00;
    mem[1901] = 8'h00;
    mem[1902] = 8'h00;
    mem[1903] = 8'h00;
    mem[1904] = 8'h00;
    mem[1905] = 8'h00;
    mem[1906] = 8'h00;
    mem[1907] = 8'h00;
    mem[1908] = 8'h00;
    mem[1909] = 8'h00;
    mem[1910] = 8'h00;
    mem[1911] = 8'h1f;
    mem[1912] = 8'h3c;
    mem[1913] = 8'h00;
    mem[1914] = 8'h00;
    mem[1915] = 8'h00;
    mem[1916] = 8'h00;
    mem[1917] = 8'h00;
    mem[1918] = 8'h00;
    mem[1919] = 8'h00;
    mem[1920] = 8'h00;
    mem[1921] = 8'h00;
    mem[1922] = 8'h00;
    mem[1923] = 8'h00;
    mem[1924] = 8'h00;
    mem[1925] = 8'h00;
    mem[1926] = 8'h00;
    mem[1927] = 8'h1e;
    mem[1928] = 8'h18;
    mem[1929] = 8'h00;
    mem[1930] = 8'h00;
    mem[1931] = 8'h00;
    mem[1932] = 8'h00;
    mem[1933] = 8'h00;
    mem[1934] = 8'h00;
    mem[1935] = 8'h00;
    mem[1936] = 8'h00;
    mem[1937] = 8'h00;
    mem[1938] = 8'h00;
    mem[1939] = 8'h00;
    mem[1940] = 8'h00;
    mem[1941] = 8'h00;
    mem[1942] = 8'h00;
    mem[1943] = 8'h1c;
    mem[1944] = 8'h0c;
    mem[1945] = 8'h00;
    mem[1946] = 8'h00;
    mem[1947] = 8'h00;
    mem[1948] = 8'h00;
    mem[1949] = 8'h00;
    mem[1950] = 8'h00;
    mem[1951] = 8'h00;
    mem[1952] = 8'h00;
    mem[1953] = 8'h00;
    mem[1954] = 8'h00;
    mem[1955] = 8'h00;
    mem[1956] = 8'h00;
    mem[1957] = 8'h00;
    mem[1958] = 8'h00;
    mem[1959] = 8'h18;
    mem[1960] = 8'h0c;
    mem[1961] = 8'h00;
    mem[1962] = 8'h00;
    mem[1963] = 8'h00;
    mem[1964] = 8'h00;
    mem[1965] = 8'h00;
    mem[1966] = 8'h00;
    mem[1967] = 8'h00;
    mem[1968] = 8'h00;
    mem[1969] = 8'h00;
    mem[1970] = 8'h00;
    mem[1971] = 8'h00;
    mem[1972] = 8'h00;
    mem[1973] = 8'h00;
    mem[1974] = 8'h00;
    mem[1975] = 8'h18;
    mem[1976] = 8'h00;
    mem[1977] = 8'h00;
    mem[1978] = 8'h00;
    mem[1979] = 8'h00;
    mem[1980] = 8'h00;
    mem[1981] = 8'h00;
    mem[1982] = 8'h00;
    mem[1983] = 8'h00;
    mem[1984] = 8'h00;
    mem[1985] = 8'h00;
    mem[1986] = 8'h00;
    mem[1987] = 8'h00;
    mem[1988] = 8'h00;
    mem[1989] = 8'h00;
    mem[1990] = 8'h00;
    mem[1991] = 8'h00;
    mem[1992] = 8'h00;
    mem[1993] = 8'h00;
    mem[1994] = 8'h00;
    mem[1995] = 8'h00;
    mem[1996] = 8'h00;
    mem[1997] = 8'h00;
    mem[1998] = 8'h00;
    mem[1999] = 8'h00;
    mem[2000] = 8'h00;
    mem[2001] = 8'h00;
    mem[2002] = 8'h00;
    mem[2003] = 8'h00;
    mem[2004] = 8'h00;
    mem[2005] = 8'h00;
    mem[2006] = 8'h00;
    mem[2007] = 8'h00;
    mem[2008] = 8'h00;
    mem[2009] = 8'h00;
    mem[2010] = 8'h00;
    mem[2011] = 8'h00;
    mem[2012] = 8'h00;
    mem[2013] = 8'h00;
    mem[2014] = 8'h00;
    mem[2015] = 8'h00;
    mem[2016] = 8'h00;
    mem[2017] = 8'h00;
    mem[2018] = 8'h00;
    mem[2019] = 8'h00;
    mem[2020] = 8'h00;
    mem[2021] = 8'h00;
    mem[2022] = 8'h00;
    mem[2023] = 8'h00;
    mem[2024] = 8'h00;
    mem[2025] = 8'h00;
    mem[2026] = 8'h00;
    mem[2027] = 8'h00;
    mem[2028] = 8'h00;
    mem[2029] = 8'h00;
    mem[2030] = 8'h00;
    mem[2031] = 8'h00;
    mem[2032] = 8'h00;
    mem[2033] = 8'h00;
    mem[2034] = 8'h00;
    mem[2035] = 8'h00;
    mem[2036] = 8'h00;
    mem[2037] = 8'h00;
    mem[2038] = 8'h00;
    mem[2039] = 8'h00;
    mem[2040] = 8'h00;
    mem[2041] = 8'h00;
    mem[2042] = 8'h00;
    mem[2043] = 8'h00;
    mem[2044] = 8'h00;
    mem[2045] = 8'h00;
    mem[2046] = 8'h00;
    mem[2047] = 8'h00;
  end

  wire [10:0] addr = {y[6:0], x[6:3]};
  assign pixel = mem[addr][x&7];

endmodule
